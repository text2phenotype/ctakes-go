aardwolves|aardwolf
abaci|abacus
aboideaux|aboideau
aboiteaux|aboiteau
abscissae|abscissa
acanthi|acanthus
acari|acarus
acciaccature|acciaccatura
acetabula|acetabulum
achaemenidae|achaemenid
achaemenides|achaemenid
aciculae|acicula
acicula|aciculum
acini|acinus
acre-feet|acre-foot
acromia|acromion
actiniae|actinia
actinozoa|actinozoan
addenda|addendum
adenocarcinomata|adenocarcinoma
adenomata|adenoma
adieux|adieu
adyta|adytum
aecia|aecium
aecidia|aecidium
aerobia|aerobium
agents-general|agent-general
aggiornamenti|aggiornamento
agnomina|agnomen
agones|agon
agorae|agora
agouties|agouti
aides-de-camp|aide-de-camp
aides-memoire|aide-memoire
aids-de-camp|aid-de-camp
alae|ala
alewives|alewife
alkalies|alkali
allodia|allodium
alluvia|alluvium
alodia|alodium
alto-relievos|alto-relievo
alto-rilievo|alto-relievo
altocumuli|altocumulus
altostrati|altostratus
alulae|alula
alumnae|alumna
alumni|alumnus
alveoli|alveolus
amanuenses|amanuensis
ambulacra|ambulacrum
amebae|ameba
amici_curiae|amicus_curiae
amnia|amnion
amniocenteses|amniocentesis
amoebae|amoeba
amoebiases|amoebiasis
amoraim|amora
amoretti|amoretto
amorini|amorino
amphiarthroses|amphiarthrosis
amphicia|amphithecium
amphimixes|amphimixis
amphioxi|amphioxus
amphisbaenae|amphisbaena
amphorae|amphora
ampullae|ampulla
amygdalae|amygdala
anabases|anabasis
anacolutha|anacoluthon
anacruses|anacrusis
anaerobia|anaerobium
anagnorises|anagnorisis
analemmata|analemma
analyses|analysis
anamneses|anamnesis
anamorphoses|anamorphosis
anastomoses|anastomosis
anatyxes|anaptyxis
ancones|ancon
ancone|ancon
androclinia|androclinium
androecia|androecium
androsphinges|androsphinx
andtheridia|antheridium
angelfishes|angelfish
angiomata|angioma
animalcula|animalculum
anlagen|anlage
annattos|anatto
annatto|anatto
annuli|annulus
antae|anta
antalkalies|antalkali
antefixa|antefix
antennae|antenna
antependia|antependium
anthelia|anthelion
anthelices|anthelix
anthemia|anthemion
antheridia|antheridium
anthodia|anthodium
anthozoa|anthozoan
anthraces|anthrax
anticlinoria|anticlinorium
antihelices|antihelix
antiheroes|antihero
antisera|antiserum
antitheses|antithesis
antitragi|antitragus
antra|antrum
anus|anus
aortae|aorta
aphelia|aphelion
aphides|aphis
apices|apex
apodoses|apodosis
apomixes|apomixis
aponeuroses|aponeurosis
apophyses|apophysis
aposiopeses|aposiopesis
apothecia|apothecium
apotheoses|apotheosis
apparatus|apparatus
appendices|appendix
appoggiature|appoggiatura
apsides|apsis
aquae|aqua
aquaria|aquarium
araglis|argali
arboreta|arboretum
arcana|arcanum
archegonia|archegonium
archerfishes|archerfish
archesporia|archesporium
archipelagoes|archipelago
arcs-boutants|arc-boutant
areolae|areola
argali|argali
argumenta|argumentum
ariette|arietta
aristae|arista
armamentaria|armamentarium
arses|arsis
artal|rotl
artel|rotl
arterioscleroses|arteriosclerosis
aruspices|aruspex
asceses|ascesis
ascidia|ascidium
asci|ascus
ascogonia|ascogonium
ashes|ash
ashkenazim|ashkenazi
aspergilla|aspergillum
aspergilli|aspergillus
aspergilloses|aspergillosis
aspersoria|aspersorium
assegais|assagai
assegai|assagai
astragali|astragalus
asyndeta|asyndeton
atheromata|atheroma
atheroscleroses|atherosclerosis
atmolyses|atmolysis
atria|atrium
attorneys-at-law|attorney-at-law
auditoria|auditorium
aurae|aura
aurar|eyrir
aurei|aureus
auriculae|auricula
aurorae|aurora
auspices|auspex
auspice|auspex
autocatalyses|autocatalysis
autochthones|autochthon
automata|automaton
autos-da-fe|auto-da-fe
avitaminoses|avitaminosis
axes|ax
axillae|axilla
axis|ax
bacchantes|bacchant
bacchante|bacchant
bacchii|bacchius
bacilli|bacillus
bacteriostases|bacteriostasis
bacula|baculum
bains-marie|bain-marie
bains_marie|bain_marie
ballistae|ballista
bambini|bambino
bandeaux|bandeau
banditti|bandit
bani|ban
banjoes|banjo
barklice|barklouse
barramundies|barramundi
bases-on-balls|base_on_balls
bases_on_balls|base_on_balls
bases|base
basidia|basidium
basileis|basileus
basis|base
bassi|basso
bastinadoes|bastinado
bateaux|bateau
batfishes|batfish
beadsmen|beadsman
beaux|beau
beches-de-mer|beche-de-mer
bedesman|beadsman
beeves|beef
behooves|behoof
bersaglieri|bersagliere
bhishties|bheesty
bhishti|bheesty
bibliothecae|bibliotheca
bicennaries|bicentenary
bicentennial|bicentenary
bijoux|bijou
bilboes|bilbo
billets-doux|billet-doux
billfishes|billfish
bimboes|bimbo
bisectrices|bisectrix
blackfeet|blackfoot
blackfishes|blackfish
blastemata|blastema
blastulae|blastula
blindfishes|blindfish
blowfishes|blowfish
bluefishes|bluefish
boarfishes|boarfish
bok|boschbok
boleti|boletus
bolivares|bolivar
bolsheviki|bolshevik
bonefishes|bonefish
bongoes|bongo
bonitoes|bonito
booklice|booklouse
bookshelves|bookshelf
boraces|borax
borborygmi|borborygmus
bordereaux|bordereau
botargoes|botargo
box-kodaks|box_kodak
boxfishes|boxfish
brachia|brachium
brainchildren|brainchild
branchiae|branchia
brants|brant
bravadoes|bravado
bravoes|bravo
bregmata|bregma
brent|brant
brethren|brother
broadcast_media|broadcast_medium
broadleaves|broadleaf
bronchi|bronchus
brothers-in-law|brother-in-law
bryozoa|bryozoan
buboes|bubo
buckoes|bucko
buckteeth|bucktooth
buffaloes|buffalo
bullae|bulla
bunde|bund
bureaux_de_change|bureau_de_change
bureaux|bureau
bursae|bursa
bushboks|boschbok
bushbok|boschbok
busses|bus
butterfishes|butterfish
byssi|byssus
cacti|cactus
caducei|caduceus
caeca|caecum
caesurae|caesura
calami|calamus
calathi|calathus
calcanei|calcaneum
calcaneus|calcaneum
calces|calx
calculi|calculus
caldaria|caldarium
calices|calix
calicoes|calico
calli|callus
calves|calf
calyces|calyx
cambia|cambium
camerae|camera
canaliculi|canaliculus
candelabra|candelabrum
candlefishes|candlefish
canthi|canthus
canulae|canula
canzoni|canzone
capita|caput
capitula|capitulum
capricci|capriccio
carabinieri|carabiniere
carbonadoes|carbonado
carcinomata|carcinoma
cargoes|cargo
carides|caryatid
carinae|carina
caroli|carolus
carpi|carpus
carpogonia|carpogonium
carryings-on|carrying-on
caryopses|caryopsis
caryopsides|caryopsis
castrati|castrato
catabases|catabasis
cataclases|cataclasis
cataloes|catalo
catalyses|catalysis
catenae|catena
catfishes|catfish
cathari|cathar
cathexes|cathexis
cattaloes|cattalo
caudices|caudex
caules|caulis
cavatine|cavatina
cavefishes|cavefish
cavetti|cavetto
cavo-rilievi|cavo-rilievo
ceca|cecum
cellae|cella
cembali|cembalo
centesimi|centesimo
centra|centrum
cephalothoraces|cephalothorax
cercariae|cercaria
cercariiae|cercaria
cerci|cercus
cerebella|cerebellum
cerebra|cerebrum
cervices|cervix
cestuses|caestus
cesurae|cesura
chadarim|cheder
chaetae|chaeta
chaises_longues|chaise_longue
chalazae|chalaza
challoth|hallah
chalutzim|chalutz
chapaties|chapati
chapatties|chapatti
chapeaux|chapeau
chasidim|chasid
chassidim|chassid
chateaux|chateau
chazanim|chazan
chedarim|cheder
chefs-d'ouvre|chef-d'ouvre
chelae|chela
chelicerae|chelicera
cherubim|cherub
chevaux-de-frise|cheval-de-frise
chiasmata|chiasma
chiasmi|chiasmus
children|child
chillies|chilli
chinese_eddoes|chinese_eddo
chitarroni|chitarrone
chlamydes|chlamys
chlamyses|chlamys
chondromata|chondroma
choragi|choragus
choriambi|choriambus
choux|chou
chromonemata|chromonema
chrysalides|chrysalis
chuvashes|chuvash
ciboria|ciborium
cicadae|cicada
cicale|cicala
cicatrices|cicatrix
ciceroni|cicerone
cicisbei|cicisbeo
cilia|cilium
cimices|cimex
cineraria|cinerarium
cingula|cingulum
cirri|cirrus
cirrocumuli|cirrocumulus
cirrostrati|cirrostratus
ciscoes|cisco
cisternae|cisterna
clani|clarino
clanos|clarino
claroes|claro
clepsydrae|clepsydra
clinandria|clinandrium
clingfishes|clingfish
clitella|clitellum
cloacae|cloaca
clostridia|clostridium
cloverleaves|cloverleaf
clypei|clypeus
coagula|coagulum
coalfishes|coalfish
cocci|coccus
coccyges|coccyx
cochleae|cochlea
codfishes|codfish
codices|codex
coelentera|coelenteron
coenuri|coenurus
cognomina|cognomen
cognosenti|cognosente
cola|colon
coleorhizae|coleorhiza
collegia|collegium
colloquia|colloquium
colluvia|colluvium
collyria|collyrium
colones|colon
colossi|colossus
columbaria|columbarium
columellae|columella
comae|coma
comatulae|comatula
comedones|comedo
comics|comic_strip
comic|comic_strip
commandoes|commando
concertanti|concertante
concerti_grossi|concerto_grosso
concertini|concertino
concerti|concerto
conchae|concha
condottieri|condottiere
condylomata|condyloma
confervae|conferva
congii|congius
conidia|conidium
conjunctivae|conjunctiva
conquistadores|conquistador
consortia|consortium
contagia|contagium
continua|continuum
contralti|contralto
conversazioni|conversazione
convolvuli|convolvulus
cooks-general|cook-general
copulae|copula
corbiculae|corbicula
coria|corium
corneae|cornea
cornua|cornu
coronae|corona
corpora_lutea|corpus_luteum
corpora_striata|corpus_striatum
corpora|corpus
corrigenda|corrigendum
cortices|cortex
cortinae|cortina
corybantes|corybant
coryphaei|coryphaeus
costae|costa
cothurni|cothurnus
courts_martial|court_martial
couteaux|couteau
cowfishes|cowfish
coxae|coxa
cramboes|crambo
crania|cranium
crases|crasis
crawfishes|crawfish
crayfishes|crayfish
credenda|credendum
crematoria|crematorium
crescendi|crescendo
cribella|cribellum
crises|crisis
crissa|crissum
cristae|crista
criteria|criterion
cruces|crux
crura|crus
crusadoes|crusado
cruzadoes|cruzado
cryings|cry
crying|cry
ctenidia|ctenidium
cubicula|cubiculum
culices|culex
culpae|culpa
culs-de-sac|cul-de-sac
culti|cultus
cumuli|cumulus
cumulonimbi|cumulonimbus
cumulostrati|cumulostratus
curiae|curia
curricula|curriculum
custodes|custos
cutes|cutis
cuticulae|cuticula
cuttlefishes|cuttlefish
cyclopes|cyclops
cycloses|cyclosis
cylices|cylix
cylikes|cylix
cymae|cyma
cymatia|cymatium
cypselae|cypsela
cysticerci|cysticercus
dadoes|dado
dagoes|dago
damselfishes|damselfish
data|datum
daughters-in-law|daughter-in-law
daymios|daimio
daymio|daimio
dealfishes|dealfish
decemviri|decemvir
decennia|decennium
deciduae|decidua
definienda|definiendum
definientia|definiens
delphinia|delphinium
denarii|denarius
dentalia|dentalium
dermatoses|dermatosis
desiderata|desideratum
desperadoes|desperado
devilfishes|devilfish
diaereses|diaeresis
diaerses|diaeresis
diagnoses|diagnosis
dialyses|dialysis
diaphyses|diaphysis
diapophyses|diapophysis
diarthroses|diarthrosis
diastalses|diastalsis
diastases|diastasis
diastemata|diastema
diathses|diathesis
diazoes|diazo
dibbukkim|dibbuk
dichasia|dichasium
dicta|dictum
didoes|dido
diereses|dieresis
dieses|diesis
differentiae|differentia
dilettanti|dilettante
diluvia|diluvium
dingoes|dingo
diplococci|diplococcus
directors-general|director-general
disci|discus
discoboli|discobolos
discobolus|discobolos
diverticula|diverticulum
divertimenti|divertimento
dive|diva
djinny|djinni
djinn|djinni
dodoes|dodo
dogfishes|dogfish
dogmata|dogma
dogteeth|dogtooth
dollarfishes|dollarfish
domatia|domatium
dominoes|domino
dormice|dormouse
dorsa|dorsum
drachmae|drachma
drawknives|drawknife
drosophilae|drosophila
drumfishes|drumfish
dryades|dryad
dui|duo
duonas|duodenum
duona|duodenum
dupondii|dupondius
duumviri|duumvir
dwarves|dwarf
dybbukkim|dybbuk
ecchymoses|ecchymosis
ecclesiae|ecclesia
ecdyses|ecdysis
echidnae|echidna
echini|echinus
echinococci|echinococcus
echoes|echo
ectozoa|ectozoan
eddoes|eddo
edemata|edema
effluvia|effluvium
eidola|eidolon
eisegeses|eisegesis
eisteddfodau|eisteddfod
elenchi|elenchus
ellipses|ellipsis
eluvia|eluvium
elves|elf
elytra|elytron
elytrum|elytron
embargoes|embargo
emboli|embolus
emphases|emphasis
emporia|emporium
enarthroses|enarthrosis
encephala|encephalon
encephalitides|encephalitis
encephalomata|encephaloma
enchiridia|enchiridion
enchondromata|enchondroma
encomia|encomium
endamebae|endameba
endamoebae|endamoeba
endocardia|endocardium
endocrania|endocranium
endometria|endometrium
endostea|endosteum
endostoses|endostosis
endothecia|endothecium
endothelia|endothelium
endotheliomata|endothelioma
endozoa|endozoan
enemata|enema
enneahedra|enneahedron
entamebae|entameba
entamoebae|entamoeba
entases|entasis
entera|enteron
entia|ens
entozoa|entozoan
entozoon|entozoan
epencephala|epencephalon
epentheses|epenthesis
epexegeses|epexegesis
ephemerae|ephemera
ephemera|ephemeron
ephemerides|ephemeris
ephori|ephor
epicalyces|epicalyx
epicanthi|epicanthus
epicardia|epicardium
epicedia|epicedium
epicleses|epiclesis
epididymides|epididymis
epigastria|epigastrium
epiglottides|epiglottis
epimysia|epimysium
epiphenomena|epiphenomenon
epiphyses|epiphysis
episterna|episternum
epithalamia|epithalamion
epithalamium|epithalamion
epithelia|epithelium
epitheliomata|epithelioma
epizoa|epizoan
epizoon|epizoan
epyllia|epyllion
equilibria|equilibrium
equiseta|equisetum
eringoes|eringo
errata|erratum
eryngoes|eryngo
esophagi|esophagus
etyma|etymon
eucalypti|eucalyptus
eupatridae|eupatrid
euripi|euripus
exanthemata|exanthema
executrices|executrix
exegeses|exegesis
exempla|exemplum
exordia|exordium
exostoses|exostosis
extrema|extremum
eyeteeth|eyetooth
fabliaux|fabliau
faciae|facia
faculae|facula
faeroese|faeroese
fallfishes|fallfish
famuli|famulus
farmers-general|farmer-general
faroese|faroese
farragoes|farrago
fasciae|fascia
fasciculi|fasciculus
fathers-in-law|father-in-law
fatsoes|fatso
faunae|fauna
feculae|fecula
fedayeen|fedayee
feet|foot
fellaheen|fellah
fellahin|fellah
felones_de_se|felo_de_se
felos_de_se|felo_de_se
femora|femur
fenestellae|fenestella
fenestrae|fenestra
feriae|feria
fermate|fermata
ferulae|ferula
festschriften|festschrift
fetiales|fetial
fezzes|fez
fiascoes|fiasco
fibrillae|fibrilla
fibromata|fibroma
fibulae|fibula
ficoes|fico
fideicommissa|fideicommissum
fieldmice|fieldmouse
figs.|fig.
filariiae|filaria
fila|filum
filefishes|filefish
fimbriae|fimbria
fishes|fish
fishwives|fishwife
fistulae|fistula
flabella|flabellum
flagella|flagellum
flagstaves|flagstaff
flambeaux|flambeau
flamines|flamen
flamingoes|flamingo
flatfeet|flatfoot
flatfishes|flatfish
fleurs-de-lis|fleur-de-lis
fleurs-de-lys|fleur-de-lys
flights_of_stairs|flight_of_stairs
flittermice|flittermouse
flocci|floccus
flocculi|flocculus
florae|flora
floreant.|floreat
florilegia|florilegium
flowers-de-luce|flower-de-luce
flyleaves|flyleaf
foci|focus
folia|folium
foramina|foramen
fora|forum
forceps|forceps
forefeet|forefoot
foreteeth|foretooth
formicaria|formicarium
formulae|formula
fornices|fornix
fortes|fortis
fossae|fossa
foveae|fovea
foveolae|foveola
fractocumuli|fractocumulus
fractostrati|fractostratus
fraena|fraenum
frauen|frau
frena|frenum
frenula|frenulum
frescoes|fresco
fricandeaux|fricandeau
fricandoes|fricando
frijoles|frijol
frogfishes|frogfish
frontes|frons
frusta|frustum
fuci|fucus
fulcra|fulcrum
fumatoria|fumatorium
fundi|fundus
fungi|fungus
funiculi|funiculus
furculae|furcula
furcula|furculum
furfures|furfur
galeae|galea
gambadoes|gambado
gametangia|gametangium
gametoecia|gametoecium
gammadia|gammadion
ganglia|ganglion
garfishes|garfish
gasses|gas
gastrulae|gastrula
gas|gas
gateaux|gateau
gazeboes|gazebo
geckoes|gecko
geese|goose
gelsemia|gelsemium
gemboks|gemsbok
gembucks|gemsbuck
gemeinschaften|gemeinschaft
gemmae|gemma
generatrices|generatrix
genera|genus
geneses|genesis
genii|genius
gentes|gens
gentlemen-at-arms|gentleman-at-arms
gentlemen-farmers|gentleman-farmer
genua|genu
genus|genus
germina|germen
gesellschaften|gesellschaft
gestalten|gestalt
ghettoes|ghetto
gingivae|gingiva
gingkoes|gingko
ginglymi|ginglymus
ginkgoes|ginkgo
gippoes|gippo
glabellae|glabella
gladioli|gladiolus
glandes|glans
gliomata|glioma
glissandi|glissando
globefishes|globefish
globigerinae|globigerina
glochidcia|glochidium
glochidia|glochidium
glomeruli|glomerulus
glossae|glossa
glottides|glottis
glutaei|glutaeus
glutei|gluteus
gnoses|gnosis
goatfishes|goatfish
goboes|gobo
godchildren|godchild
goes|go
goings-over|going-over
goldfishes|goldfish
gomphoses|gomphosis
gonia|gonion
gonidia|gonidium
gonococci|gonococcus
goodwives|goodwife
goosefishes|goosefish
gorgoneia|gorgoneion
gospopoda|gospodin
governors_general|governor_general
goyim|goy
gps|gps
grafen|graf
graffiti|graffito
grandchildren|grandchild
grants-in-aid|grant-in-aid
granulomata|granuloma
gravamina|gravamen
grig-gris|gris-gris
groszy|grosz
grottoes|grotto
guilders|guilde
guilder|guilde
guitarfishes|guitarfish
gummata|gumma
gurnards|gurnar
gurnard|gurnar
guttae|gutta
gymnasia|gymnasium
gynaecea|gynaeceum
gynaecia|gynaecium
gynecea|gynecium
gynecia|gynecium
gynoecea|gynoecium
gynoecia|gynoecium
gyri|gyrus
hadarim|heder
hadjes|hadj
haematolyses|haematolysis
haematomata|haematoma
haematozoa|haematozoon
haemodialyses|haemodialysis
haemolyses|haemolysis
haemoptyses|haemoptysis
haeredes|haeres
haftaroth|haftarah
hagfishes|hagfish
haggadah|haggada
haggadas|haggada
haggadoth|haggada
hajjes|hajj
haleru|haler
halfpence|halfpenny
halloth|hallah
hallot|hallah
halluces|hallux
haloes|halo
halteres|halter
haltere|halter
halves|half
hamuli|hamulus
hangers-on|hanger-on
haphtaroth|haphtarah
haredim|haredi
haruspices|haruspex
hasidim|hasid
hassidim|hassid
haustella|haustellum
haustoria|haustorium
hazzanim|hazzan
hectocotyli|hectocotylus
heirs-at-law|heir-at-law
heldentenore|heldentenor
helices|helix
heliozoa|heliozoan
hematolyses|hematolysis
hematomata|hematoma
hematozoa|hematozoon
hemelytra|hemelytron
hemielytra|hemielytron
hemodialyses|hemodialysis
hemolyses|hemolysis
hemoptyses|hemoptysis
hendecahedra|hendecahedron
hens-and-chickens|hen-and-chickens
heraclidae|heraclid
heraklidae|heraklid
herbaria|herbarium
hermae|herm
hermai|herma
herma|herm
herniae|hernia
heroes|hero
herren|herr
hetaerae|hetaera
hetairai|hetaira
hibernacula|hibernaculum
hieracosphinges|hieracosphinx
hila|hilum
hili|hilus
himatia|himation
hippocampi|hippocampus
hippopotami|hippopotamus
his|his
hoboes|hobo
hogfishes|hogfish
homunculi|homunculus
honoraria|honorarium
hooves|hoof
horologia|horologium
houses_of_cards|house_of_cards
housewives|housewife
humeri|humerus
hydrae|hydra
hydromedusae|hydromedusa
hydrozoa|hydrozoan
hymenoptera|hymenopteran
hynia|hymenium
hyniums|hymenium
hypanthia|hypanthium
hyperostoses|hyperostosis
hyphae|hypha
hypnoses|hypnosis
hypochondria|hypochondrium
hypogastria|hypogastrium
hypogea|hypogeum
hypophyses|hypophysis
hypostases|hypostasis
hypothalami|hypothalamus
hypotheses|hypothesis
hyraces|hyrax
iambi|iamb
ibices|ibex
ibo|igbo
ichthyosauri|ichthyosaurus
ichthyosauruses|ichthyosaur
ichthyosaurus|ichthyosaur
iconostases|iconostas
iconostasis|iconostas
icosahedra|icosahedron
ideata|ideatum
igorrorote|igorrote
ilia|ilium
imagines|imago
imagoes|imago
imperia|imperium
impies|impi
incubi|incubus
incudes|incus
indices|index
indigoes|indigo
indumenta|indumentum
indusia|indusium
infundibula|infundibulum
ingushes|ingush
innuendoes|innuendo
inocula|inoculum
inquisitors-general|inquisitor-general
insectaria|insectarium
insulae|insula
intagli|intaglio
interleaves|interleaf
intermezzi|intermezzo
interreges|interrex
interregna|interregnum
intimae|intima
involucella|involucellum
involucra|involucrum
irides|iris
irs|irs
ischia|ischium
isthmi|isthmus
is|is
jackeroos|jackaroo
jackeroo|jackaroo
jackfishes|jackfish
jackknives|jackknife
jacks-in-the-box|jack-in-the-box
jambeaux|jambeau
jellyfishes|jellyfish
jewelfishes|jewelfish
jewfishes|jewfish
jingoes|jingo
jinn|jinni
joes|jo
joe|jo
judge_advocates_general|judge_advocate_general
jura|jus
kaddishim|kaddish
kalmucks|kalmuc
kalmuck|kalmuc
katabases|katabasis
keeshonden|keeshond
kibbutzim|kibbutz
killifishes|killifish
kingfishes|kingfish
kings-of-arms|king-of-arms
knights_bachelors|knight_bachelor
knights_bachelor|knight_bachelor
knights_templars|knight_templar
knights_templar|knight_templar
knives|knife
kohlrabies|kohlrabi
kronen|krone
kroner|krone
kronur|krona
krooni|kroon
kylikes|kylix
labara|labarum
labella|labellum
labia|labium
labra|labrum
lactobacilli|lactobacillus
lacunae|lacuna
lacunaria|lacunar
ladies-in-waiting|lady-in-waiting
lamellae|lamella
lamiae|lamia
laminae|lamina
lapilli|lapillus
lapithae|lapith
larvae|larva
larynges|larynx
lassoes|lasso
latices|latex
latifundia|latifundium
lati|lat
latu|lat
lavaboes|lavabo
leaves|leaf
leave|leaf
lecythi|lecythus
leges|lex
lei|leu
lemmata|lemma
lemnisci|lemniscus
lenes|lenis
lentigines|lentigo
leonides|leonid
lepidoptera|lepidopteran
leprosaria|leprosarium
lepta|lepton
leptocephali|leptocephalus
leucocytozoa|leucocytozoan
leva|lev
librae|libra
libretti|libretto
lice|louse
lieder|lied
ligulae|ligula
limbi|limbus
limina|limen
limites|limes
limuli|limulus
lingoes|lingo
linguae_francae|lingua_franca
linguae|lingua
lionfishes|lionfish
lipomata|lipoma
lire|lira
liriodendra|liriodendron
lisente|sente
listente|sente
litai|lit
litas|lit
litu|litas
lives|life
lixivia|lixivium
loaves|loaf
loci|locus
loculi|loculus
loggie|loggia
logia|logion
lomenta|lomentum
longobardi|longobard
loricae|lorica
loups-garous|loup-garou
luba|luba
lubritoria|lubritorium
lumbus|lumbi
lumina|lumen
lumpfishes|lumpfish
lungfishes|lungfish
lunulae|lunula
lures|lur
lure|lur
lustra|lustre
lyings-in|lying-in
lymphangitides|lymphangitis
lymphomata|lymphoma
lymphopoieses|lymphopoiesis
lyses|lysis
lyttae|lytta
maare|maar
macaronies|macaroni
maccaronies|maccaroni
machzorim|machzor
macronuclei|macronucleus
macrosporangia|macrosporangium
maculae|macula
madornos|madrono
maestri|maestro
mafiosi|mafioso
magi|magus
magmata|magma
magnificoes|magnifico
mahzorim|mahzor
major-axes|major_axis
major_axes|major_axis
makuta|likuta
mallei|malleus
malleoli|malleolus
maloti|loti
mamillae|mamilla
mammae|mamma
mammillae|mammilla
mandingoes|mandingo
mangoes|mango
manifestoes|manifesto
manteaux|manteau
mantes|mantis
manubria|manubrium
marchese|marchesa
marchesi|marchese
maremme|maremma
markkaa|markka
marsupia|marsupium
marvels-of-peru|marvel-of-peru
mass_media|mass_medium
masses|mass
masse|mass
masters-at-arms|master-at-arms
matrices|matrix
matzoth|matzo
mausolea|mausoleum
maxillae|maxilla
maxima|maximum
mediae|media
mediastina|mediastinum
media|medium
medullae_oblongatae|medulla_oblongata
medullae|medulla
medusae|medusa
megara|megaron
megasporangia|megasporangium
megilloth|megillah
meioses|meiosis
melanomata|melanoma
melismata|melisma
mementoes|memento
memoranda|memorandum
men-at-arms|man-at-arms
men-o'-war|man-of-war
men-of-war|man-of-war
men_of_letters|man_of_letters
menisci|meniscus
menservants|manservant
menstrua|menstruum
men|man
mesdames|madame
mesdemoiselles|mademoiselle
mesentera|mesenteron
mesothoraces|mesothorax
messeigneurs|monseigneur
messieurs|monsieur
mestizoes|mestizo
metacarpi|metacarpus
metamorphoses|metamorphosis
metanephroi|metanephros
metastases|metastasis
metatarsi|metatarsus
metatheses|metathesis
metathoraces|metathorax
metazoa|metazoan
metempsychoses|metempsychosis
metencephala|metencephalon
mezuzoth|mezuzah
miasmata|miasma
mice|mouse
microanalyses|microanalysis
micrococci|micrococcus
micronuclei|micronucleus
microsporangia|microsporangium
midrashim|midrash
midwives|midwife
milia|milium
milieux|milieu
militated_against|militate_against
milkfishes|milkfish
millennia|millennium
minae|mina
minima|minimum
ministeria|ministerium
minutiae|minutia
minyanim|minyan
mioses|miosis
miracidia|miracidium
miri|mir
mishnah|mishna
mishnayoth|mishna
mitochondria|mitochondrion
mitzvoth|mitzvah
modioli|modiolus
moduli|modulus
momenta|momentum
moments_of_truth|moment_of_truth
momi|momus
monades|monad
monas|monad
monkfishes|monkfish
monochasia|monochasium
monopodia|monopodium
monoptera|monopteron
monopteroi|monopteros
monsignori|monsignor
monts-de-piete|mont-de-piete
mooncalves|mooncalf
moonfishes|moonfish
morae|mora
moratoria|moratorium
morceaux|morceau
morescoes|moresco
moriscoes|morisco
morphallaxes|morphallaxis
morphoses|morphosis
morses|morse
mors|morse
morulae|morula
mosasauri|mosasaurus
moshavim|moshav
moslims|moslem
moslim|moslem
mosquitoes|mosquito
mothers-in-law|mother-in-law
mothers_superior|mother_superior
mottoes|motto
movers_and_shakers|mover_and_shaker
mucosae|mucosa
mucrones|mucro
mudejares|mudejar
mudfishes|mudfish
mulattoes|mulatto
multiparae|multipara
murices|murex
muskallunge|muskellunge
mycelia|mycelium
mycetomata|mycetoma
mycobacteria|mycobacterium
mycorrhizae|mycorrhiza
myelencephala|myelencephalon
myiases|myiasis
myocardia|myocardium
myofibrillae|myofibrilla
myomata|myoma
myoses|myosis
myrmidones|myrmidon
mythoi|mythos
myxomata|myxoma
naevi|naevus
naiades|naiad
naoi|naos
narcissi|narcissus
nares|naris
nasopharynges|nasopharynx
natatoria|natatorium
naumachiae|naumachia
nauplii|nauplius
nautili|nautilus
navahoes|navaho
navajoes|navajo
nebulae|nebula
necropoleis|necropolis
needlefishes|needlefish
negrilloes|negrillo
negritoes|negrito
negroes|negro
nemeses|nemesis
nephridia|nephridium
nereides|nereid
neurohypophyses|neurohypophysis
neuromata|neuroma
neuroptera|neuropteron
neuroses|neurosis
nevi|nevus
nibelungen|nibelung
nidi|nidus
nielli|niello
nilgai|nilgai
nimbi|nimbus
nimbostrati|nimbostratus
noctilucae|noctiluca
nodi|nodus
noes|no
nomina|nomen
nota|notum
noumena|noumenon
novae|nova
novelle|novella
novenae|novena
nubeculae|nubecula
nucelli|nucellus
nuchae|nucha
nuclei|nucleus
nucleoli|nucleolus
nulliparae|nullipara
numbfishes|numbfish
numina|numen
nymphae|nympha
oarfishes|oarfish
oases|oasis
obeli|obelus
objets_d'art|objet_d'art
obligati|obligato
oboli|obolus
occipita|occiput
oceanaria|oceanarium
oceanides|oceanid
ocelli|ocellus
ochreae|ochrea
ocreae|ochrea
ocrea|ochrea
octahedra|octahedron
octopi|octopus
oculi|oculus
odea|odeum
oedemata|edema
oedema|edema
oesophagi|esophagus
oesophagus|esophagus
oldwives|oldwife
olea|oleum
omasa|omasum
omayyades|omayyad
omenta|omentum
ommatidia|ommatidium
ommiades|ommiad
onagri|onager
oogonia|oogonium
oothecae|ootheca
operas_seria|opera_seria
opercula|operculum
optic_axes|optic_axis
optima|optimum
ora|os
organa|organon
organums|organa
organum|organa
orthoptera|orthopteron
osar|os
oscula|osculum
ossa|os
osteomata|osteoma
ostia|ostium
ottomans|othman
ottoman|othman
ova|ovum
ovoli|ovolo
ovotestes|ovotestis
oxen|ox
oxymora|oxymoron
paddlefishes|paddlefish
paise|paisa
paleae|palea
palestrae|palestra
palingeneses|palingenesis
pallia|pallium
palmettoes|palmetto
palpi|palpus
pancratia|pancratium
panettoni|panettone
paparazzi|paparazzo
paperknives|paperknife
papillae|papilla
papillomata|papilloma
pappi|pappus
papulae|papula
papyri|papyrus
parabases|parabasis
paraleipses|paraleipsis
paralipsis|paraleipsis
paralyses|paralysis
paramecia|paramecium
paramenta|parament
paraphyses|paraphysis
parapodia|parapodium
parapraxes|parapraxis
paraselenae|paraselene
parashoth|parashah
parasyntheta|parasyntheton
parazoa|parazoan
parentheses|parenthesis
parerga|parergon
parhelia|parhelion
parietes|paries
paris-mutuels|pari-mutuel
parrotfishes|parrotfish
parulides|parulis
pasos_dobles|paso_doble
passers-by|passer-by
pastorali|pastorale
patagia|patagium
patellae|patella
patinae|patina
patresfamilias|paterfamilias
pease|pea
peccadilloes|peccadillo
pectines|pecten
pedaloes|pedalo
pedes|pes
pekingese|pekinese
pelves|pelvis
pence|penny
penes|penis
penetralium|penetralia
penicillia|penicillium
penknives|penknife
pennae|penna
pennia|penni
pentahedra|pentahedron
pentimenti|pentimento
penumbrae|penumbra
pepla|peplum
pericardia|pericardium
perichondria|perichondrium
pericrania|pericranium
peridia|peridium
perigonia|perigonium
perihelia|perihelion
perinea|perineum
perinephria|perinephrium
perionychia|perionychium
periostea|periosteum
periphrases|periphrasis
peristalses|peristalsis
perithecia|perithecium
peritonea|peritoneum
personae|persona
petechiae|petechia
pfennige|pfennig
phalanges|phalange
phalanx|phalange
phalli|phallus
pharynges|pharynx
phenomena|phenomenon
phi-phenomena|phi-phenomenon
philodendra|philodendron
phlyctenae|phlyctaena
phlyctena|phlyctaena
phylae|phyle
phyla|phylum
phyllotaxes|phyllotaxis
phylloxerae|phylloxera
phylogeneses|phylogenesis
pieds-a-terre|pied-a-terre
pigfishes|pigfish
pilea|pileum
pilei|pileus
pineta|pinetum
pinfishes|pinfish
pinkoes|pinko
pinnae|pinna
pinnulae|pinnula
pipefishes|pipefish
pirogi|pirog
piscinae|piscina
pithecanthropi|pithecanthropus
pithoi|pithos
placeboes|placebo
placentae|placenta
planetaria|planetarium
planulae|planula
plasmodesmata|plasmodesma
plasmodia|plasmodium
plateaux|plateau
plectra|plectron
plectrum|plectron
plena|plenum
pleurae|pleura
pleura|pleuron
plicae|plica
ploughmen|ploughman
plowman|ploughman
pneumobacilli|pneumobacillus
pneumococci|pneumococcus
pocketknives|pocketknife
podetia|podetium
podia|podium
poleis|polis
pollices|pollex
pollinia|pollinium
polychasia|polychasium
polyhedra|polyhedron
polyparia|polyparium
polypi|polypus
polyzoaria|polyzoarium
polyzoa|polyzoan
pontes|pons
pontifices|pontifex
portamenti|portamento
porticoes|portico
portmanteaux|portmanteau
postliminia|postliminium
potatoes|potato
praenomina|praenomen
praxes|praxis
predelle|predella
premaxillae|premaxilla
prenomina|prenomen
prese|presa
primigravidae|primigravida
primiparae|primipara
primi|primo
primordia|primordium
principia|principium
proboscides|proboscis
proces-verbaux|proces-verbal
proglottides|proglottid
proglottis|proglottid
prognoses|prognosis
prolegomena|prolegomenon
prolepses|prolepsis
promycelia|promycelium
pronephra|pronephros
pronephroi|pronephros
pronuclei|pronucleus
propositi|propositus
proptoses|proptosis
propylaea|propylaeum
propyla|propylon
proscenia|proscenium
prosencephala|prosencephalon
prostheses|prosthesis
prostomia|prostomium
protases|protasis
prothalamia|prothalamion
prothalamium|prothalamion
prothallia|prothallium
prothalli|prothallus
prothoraces|prothorax
protonemata|protonema
protozoa|protozoan
proventriculi|proventriculus
provisoes|proviso
prytanea|prytaneum
psalteria|psalterium
pseudopodia|pseudopodium
psychoneuroses|psychoneurosis
psychoses|psychosis
pterygia|pterygium
pterylae|pteryla
ptoses|ptosis
pubes|pubis
pudenda|pudendum
puli|pul
pulvilli|pulvillus
pulvini|pulvinus
punchinelloes|punchinello
pupae|pupa
puparia|puparium
putamina|putamen
putti|putto
pycnidia|pycnidium
pygidia|pygidium
pylori|pylorus
pyxides|pyxis
pyxidia|pyxidium
qaddishim|qaddish
quadrennia|quadrennium
quadrigae|quadriga
qualia|quale
quanta|quantum
quarterstaves|quarterstaff
quezales|quezal
quinquennia|quinquennium
quizzes|quiz
rabatos|rabato
rabbitfishes|rabbitfish
rachides|rhachis
radices|radix
radii|radius
radulae|radula
ramenta|ramentum
rami|ramus
ranulae|ranula
ranunculi|ranunculus
raphae|raphe
raphides|raphide
raphis|raphide
ratfishes|ratfish
reales|real
rearmice|rearmouse
rebato|rabato
recta|rectum
recti|rectus
rectrices|rectrix
redfishes|redfish
rediae|redia
referenda|referendum
refugia|refugium
reguli|regulus
reis|real
relata|relatum
remiges|remex
reremice|rearmouse
reremouse|rearmouse
reseaux|reseau
residua|residuum
responsa|responsum
retiarii|retiarius
retia|rete
reticula|reticulum
retinacula|retinaculum
retinae|retina
rhabdomyomata|rhabdomyoma
rhachides|rhachis
rhachises|rachis
rhachis|rachis
rhinencephala|rhinencephalon
rhizobia|rhizobium
rhombi|rhombus
rhonchi|rhonchus
rhyta|rhyton
ribbonfishes|ribbonfish
ricercacari|ricercare
ricercari|ricercare
rickettsiae|rickettsia
rilievi|rilievo
rimae|rima
robes-de-chambre|robe-de-chambre
rockfishes|rockfish
romans-fleuves|roman-fleuve
roma|rom
rondeaux|rondeau
rosaria|rosarium
rosefishes|rosefish
rostella|rostellum
rostra|rostrum
rouleaux|rouleau
rugae|ruga
rumina|rumen
runners-up|runner-up
sacraria|sacrarium
sacra|sacrum
saguaros|saguaro
sahuaro|saguaro
sailfishes|sailfish
salespeople|salesperson
salmonellae|salmonella
salpae|salpa
salpinges|salpinx
saltarelli|saltarello
salvoes|salvo
sancta|sanctum
sanitaria|sanitarium
santimi|santims
saphenae|saphena
sarcophagi|sarcophagus
sartorii|sartorius
sassanidae|sassanid
sawfishes|sawfish
scaldfishes|scaldfish
scaleni|scalenus
scapulae|scapula
scarabaei|scarabaeus
scarves|scarf
schatchonim|schatchen
schemata|schema
scherzandi|scherzando
scherzi|scherzo
schmoes|schmo
scholia|scholium
schuln|schul
schutzstaffeln|schutzstaffel
scirrhi|scirrhus
scleromata|scleroma
scleroses|sclerosis
sclerotia|sclerotium
scoleces|scolex
scolices|scolex
scopulae|scopula
scoriae|scoria
scotomata|scotoma
scriptoria|scriptorium
scrota|scrotum
scudi|scudo
scuta|scutum
scutella|scutellum
scyphistomae|scyphistoma
scyphi|scyphus
scyphozoa|scyphozoan
secondi|secondo
secretaries-general|secretary-general
segni|segno
seleucidae|seleucid
selves|self
senores|senor
sensilla|sensillum
senti|sent
senussis|senusi
senussi|senusi
separatrices|separatrix
sephardim|sephardi
septaria|septarium
septa|septum
septennia|septennium
sequelae|sequela
sequestra|sequestrum
seraphim|seraph
sera|serum
sestertia|sestertium
setae|seta
sgraffiti|sgraffito
shabbasim|shabbas
shabbatim|shabbat
shackoes|shacko
shadchanim|shadchan
shadchans|schatchen
shadchan|schatchen
shakoes|shako
shammes|shammas
shammosim|shammas
sheatfishes|sheatfish
sheaves|sheaf
shellfishes|shellfish
shelves|shelf
shinleaves|shinleaf
shittim|shittah
shmoes|shmo
shofroth|shofar
shophar|shofar
shophroth|shophar
shrewmice|shrewmouse
shuln|shul
siddurim|siddur
sigloi|siglos
signore|signior
signorine|signorina
signori|signior
siliquae|siliqua
silvae|silva
silverfishes|silverfish
simulacra|simulacrum
sincipita|sinciput
sinfonie|sinfonia
sisters-in-law|sister-in-law
sistra|sistrum
situlae|situla
smalti|smalto
snaggleteeth|snaggletooth
snailfishes|snailfish
snipefishes|snipefish
socmen|socman
sokeman|socman
solaria|solarium
solatia|solatium
sola|solum
soldi|soldo
soles|sol
sole|sol
solfeggi|solfeggio
solidi|solidus
soli|solo
somata|soma
sons-in-law|son-in-law
soprani|soprano
sordini|sordino
sori|sorus
soroses|sorosis
sovkhozy|sovkhoz
spadefishes|spadefish
spadices|spadix
spearfishes|spearfish
spectra|spectrum
specula|speculum
spermatia|spermatium
spermatogonia|spermatogonium
spermatozoa|spermatozoon
spermogonia|spermogonium
sphinges|sphinx
spicae|spica
spicula|spiculum
spirilla|spirillum
splayfeet|splayfoot
splenii|splenius
sporangia|sporangium
sporogonia|sporogonium
sporozoa|sporozoan
springhase|springhaas
spumoni|spumone
sputa|sputum
squamae|squama
squashes|squash
squillae|squilla
squirrelfishes|squirrelfish
squizzes|squiz
stadia|stadium
stamina|stamen
staminodia|staminodium
stapedes|stapes
staphylococci|staphylococcus
staretsy|starets
starfishes|starfish
startsy|starets
stelae|stele
stemmata|stemma
stenoses|stenosis
stepchildren|stepchild
sterna|sternum
stigmata|stigma
stimuli|stimulus
stipites|stipes
stirpes|stirps
stoae|stoa
stockfishes|stockfish
stomata|stoma
stomodaea|stomodaeum
stomodea|stomodeum
stonefishes|stonefish
stotinki|stotinka
stotkini|stotinka
strappadoes|strappado
strata|stratum
strati|stratus
stratocumuli|stratocumulus
street_children|street_child
streptococci|streptococcus
stretti|stretto
striae|stria
strobili|strobilus
stromata|stroma
strumae|struma
stuccoes|stucco
styli|stylus
stylopes|stylops
stylopodia|stylopodium
subcortices|subcortex
subdeliria|subdelirium
subgenera|subgenus
subindices|subindex
submucosae|submucosa
subphyla|subphylum
substrasta|substratum
succedanea|succedaneum
succubi|succubus
suckerfishes|suckerfish
suckfishes|suckfish
sudaria|sudarium
sudatoria|sudatorium
sulci|sulcus
summae|summa
sunfishes|sunfish
supercargoes|supercargo
superheroes|superhero
supernovae|supernova
superstrata|superstratum
surgeonfishes|surgeonfish
swamies|swami
sweetiewives|sweetiewife
swellfishes|swellfish
swordfishes|swordfish
syconia|syconium
syllabi|syllabus
syllepses|syllepsis
symphyses|symphysis
sympodia|sympodium
symposia|symposium
synapses|synapsis
synarthroses|synarthrosis
synclinoria|synclinorium
syncytia|syncytium
syndesmoses|syndesmosis
synopses|synopsis
syntagmata|syntagma
syntheses|synthesis
syphilomata|syphiloma
syringes|syrinx
syssarcoses|syssarcosis
tableaux|tableau
taeniae|taenia
tali|talus
tallaisim|tallith
tallithes|tallith
tallitoth|tallith
tapeta|tapetum
tarantulae|tarantula
tarsi|tarsus
tarsometatarsi|tarsometatarsus
taxa|taxon
taxes|tax
taxies|taxi
taxis|tax
tectrices|tectrix
teeth|tooth
tegmina|tegmen
telae|tela
telamones|telamon
telangiectases|telangiectasia
telangiectasis|telangiectasia
telia|telium
tempi|tempo
tenacula|tenaculum
tenderfeet|tenderfoot
teniae|tenia
tenia|taenia
tenues|tenuis
teraphim|teraph
terata|teras
teredines|teredo
terga|tergum
termini|terminus
terraria|terrarium
terzetti|terzetto
tesserae|tessera
testae|testa
testes|testis
testudines|testudo
tetrahedra|tetrahedron
tetraskelia|tetraskelion
thalamencephala|thalamencephalon
thalami|thalamus
thalli|thallus
theatres-in-the-round|theatre-in-the-round
thecae|theca
therses|thyrse
thesauri|thesaurus
theses|thesis
thickleaves|thickleaf
thieves|thief
tholoi|tholos
thoraces|thorax
thrombi|thrombus
thymi|thymus
thyrsi|thyrsus
tibiae|tibia
tilefishes|tilefish
tintinnabula|tintinnabulum
titmice|titmouse
toadfishes|toadfish
tobaccoes|tobacco
tomatoes|tomato
tomenta|tomentum
tondi|tondo
tonneaux|tonneau
tophi|tophus
topoi|topos
tori|torus
tornadoes|tornado
torpedoes|torpedo
torsi|torso
touracos|touraco
trabeculae|trabecula
tracheae|trachea
traditores|traditor
tragi|tragus
trapezia|trapezium
trapezohedra|trapezohedron
traumata|trauma
treponemata|treponema
trichinae|trichina
triclinia|triclinium
triennia|triennium
triforia|triforium
triggerfishes|triggerfish
trihedra|trihedron
triskelia|triskelion
trisoctahedra|trisoctahedron
triumviri|triumvir
trivia|trivium
trochleae|trochlea
tropaeola|tropaeolum
trous-de-loup|trou-de-loup
trousseaux|trousseau
trunkfishes|trunkfish
trymata|tryma
tubae|tuba
turaco|touraco
turves|turf
tympana|tympanum
tyros|tiro
tyro|tiro
ubermenschen|ubermensch
uglies|ugli
uigurs|uighur
ulnae|ulna
ultimata|ultimatum
umbilici|umbilicus
umbones|umbo
umbrae|umbra
uncidia|uredium
unci|uncus
uredines|uredo
uredinia|uredinium
uredosori|uredosorus
urethrae|urethra
urinalyses|urinalysis
uteri|uterus
utriculi|utriculus
uvulae|uvula
vacua|vacuum
vaginae|vagina
vagi|vagus
vagus|vagus
valleculae|vallecula
vaporetti|vaporetto
varices|varix
vasa|vas
vascula|vasculum
velamina|velamen
velaria|velarium
vela|velum
venae_cavae|vena_cava
venae|vena
ventriculi|ventriculus
vermes|vermis
verrucae|verruca
vertebrae|vertebra
vertices|vertex
vertigines|vertigo
vertigoes|vertigo
vesicae|vesica
vetoes|veto
vexilla|vexillum
viatica|viaticum
viatores|viator
vibracula|vibraculum
vibrissae|vibrissa
vice-chairman|vice-chairman
villi|villus
vimina|vimen
vincula|vinculum
viragoes|virago
vires|vis
virtuosi|virtuoso
vitae|vita
vitelli|vitellus
vittae|vitta
vivaria|vivarium
voces|vox
volcanoes|volcano
volkslieder|volkslied
volte|volta
volvae|volva
vorticellae|vorticella
vortices|vortex
vulvae|vulva
wagons-lits|wagon-lit
wahhabis|wahabi
wahhabi|wahabi
wanderjahre|wanderjahr
weakfishes|weakfish
werewolves|werewolf
wharves|wharf
whippers-in|whipper-in
whitefishes|whitefish
wives|wife
wolffishes|wolffish
wolves|wolf
woodlice|woodlouse
wreckfishes|wreckfish
wunderkinder|wunderkind
xiphisterna|xiphisternum
yeshivahs|yeshiva
yeshivoth|yeshiva
yogin|yogi
yourselves|yourself
zamindaris|zamindari
zecchini|zecchino
zemindari|zamindari
zeroes|zero
zoaeae|zoaea
zoa|zoon
zoeae|zoea
zoeas|zoaea
zoea|zoaea
zoonoses|zoonosis
zoosporangia|zoosporangium