s|
ies|y
es|e
es|
ed|e
ed|
ing|e
ing|