s|
ses|s
xes|x
zes|z
ches|ch
shes|sh
men|man
ies|y