best|well
better|well
deeper|deeply
farther|far
further|far
harder|hard
hardest|hard