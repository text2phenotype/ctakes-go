'nt_RB|not
n't_RB|not
'd_MD|would
'll_MD|will