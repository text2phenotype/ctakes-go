acer|acer
after|after
airier|airy
airiest|airy
all-arounder|all-arounder
angrier|angry
angriest|angry
archer|archer
artier|arty
artiest|arty
ashier|ashy
ashiest|ashy
assaulter|assaulter
attacker|attacker
backer|backer
baggier|baggy
baggiest|baggy
balkier|balky
balkiest|balky
balmier|balmy
balmiest|balmy
bandier|bandy
bandiest|bandy
bargainer|bargainer
barmier|barmy
barmiest|barmy
battier|batty
battiest|batty
baulkier|baulky
baulkiest|baulky
bawdier|bawdy
bawdiest|bawdy
bayer|bayer
beadier|beady
beadiest|beady
beastlier|beastly
beastliest|beastly
beater|beater
beefier|beefy
beefiest|beefy
beerier|beery
beeriest|beery
bendier|bendy
bendiest|bendy
best|good
better|good
bigger|big
biggest|big
bitchier|bitchy
bitchiest|bitchy
biter|biter
bittier|bitty
bittiest|bitty
blearier|bleary
bleariest|bleary
bloodier|bloody
bloodiest|bloody
bloodthirstier|bloodthirsty
bloodthirstiest|bloodthirsty
blowier|blowy
blowiest|blowy
blowsier|blowsy
blowsiest|blowsy
blowzier|blowzy
blowziest|blowzy
bluer|blue
bluest|blue
boner|boner
bonier|bony
boniest|bony
bonnier|bonny
bonniest|bonny
boozier|boozy
booziest|boozy
boskier|bosky
boskiest|bosky
bossier|bossy
bossiest|bossy
botchier|botchy
botchiest|botchy
bother|bother
bouncier|bouncy
bounciest|bouncy
bounder|bounder
bower|bower
brainier|brainy
brainiest|brainy
brashier|brashy
brashiest|brashy
brassier|brassy
brassiest|brassy
brawnier|brawny
brawniest|brawny
breathier|breathy
breathiest|breathy
breezier|breezy
breeziest|breezy
brinier|briny
briniest|briny
britisher|britisher
broadcaster|broadcaster
brooder|brooder
broodier|broody
broodiest|broody
bubblier|bubbly
bubbliest|bubbly
buggier|buggy
buggiest|buggy
bulkier|bulky
bulkiest|bulky
bumpier|bumpy
bumpiest|bumpy
bunchier|bunchy
bunchiest|bunchy
burlier|burly
burliest|burly
burrier|burry
burriest|burry
burster|burster
bushier|bushy
bushiest|bushy
busier|busy
busiest|busy
buster|buster
bustier|busty
bustiest|busty
cagier|cagey
cagiest|cagey
camper|camper
cannier|canny
canniest|canny
canter|canter
cantier|canty
cantiest|canty
caster|caster
catchier|catchy
catchiest|catchy
cattier|catty
cattiest|catty
cer|cer
chancier|chancy
chanciest|chancy
charier|chary
chariest|chary
chattier|chatty
chattiest|chatty
cheekier|cheeky
cheekiest|cheeky
cheerier|cheery
cheeriest|cheery
cheesier|cheesy
cheesiest|cheesy
chestier|chesty
chestiest|chesty
chewier|chewy
chewiest|chewy
chillier|chilly
chilliest|chilly
chintzier|chintzy
chintziest|chintzy
chippier|chippy
chippiest|chippy
choosier|choosy
choosiest|choosy
choppier|choppy
choppiest|choppy
chubbier|chubby
chubbiest|chubby
chuffier|chuffy
chuffiest|chuffy
chummier|chummy
chummiest|chummy
chunkier|chunky
chunkiest|chunky
churchier|churchy
churchiest|churchy
clammier|clammy
clammiest|clammy
classier|classy
classiest|classy
cleanlier|cleanly
cleanliest|cleanly
clerklier|clerkly
clerkliest|clerkly
cloudier|cloudy
cloudiest|cloudy
clubbier|clubby
clubbiest|clubby
clumsier|clumsy
clumsiest|clumsy
cockier|cocky
cockiest|cocky
coder|coder
collier|colly
colliest|colly
comelier|comely
comeliest|comely
comfier|comfy
comfiest|comfy
cornier|corny
corniest|corny
cosier|cosy
cosiest|cosy
costlier|costly
costliest|costly
costumer|costumer
counterfeiter|counterfeiter
courtlier|courtly
courtliest|courtly
cozier|cozy
coziest|cozy
crabbier|crabby
crabbiest|crabby
cracker|cracker
craftier|crafty
craftiest|crafty
craggier|craggy
craggiest|craggy
crankier|cranky
crankiest|cranky
crasher|crasher
crawlier|crawly
crawliest|crawly
crazier|crazy
craziest|crazy
creamer|creamer
creamier|creamy
creamiest|creamy
creepier|creepy
creepiest|creepy
crispier|crispy
crispiest|crispy
crumbier|crumby
crumbiest|crumby
crumblier|crumbly
crumbliest|crumbly
crummier|crummy
crummiest|crummy
crustier|crusty
crustiest|crusty
curlier|curly
curliest|curly
customer|customer
cuter|cute
daffier|daffy
daffiest|daffy
daintier|dainty
daintiest|dainty
dandier|dandy
dandiest|dandy
deadlier|deadly
deadliest|deadly
dealer|dealer
deserter|deserter
dewier|dewy
dewiest|dewy
dicier|dicey
diciest|dicey
dimer|dimer
dimmer|dim
dimmest|dim
dingier|dingy
dingiest|dingy
dinkier|dinky
dinkiest|dinky
dippier|dippy
dippiest|dippy
dirtier|dirty
dirtiest|dirty
dishier|dishy
dishiest|dishy
dizzier|dizzy
dizziest|dizzy
dodgier|dodgy
dodgiest|dodgy
dopier|dopey
dopiest|dopey
dottier|dotty
dottiest|dotty
doughier|doughy
doughiest|doughy
doughtier|doughty
doughtiest|doughty
dowdier|dowdy
dowdiest|dowdy
dowier|dowie
dowiest|dowie
downer|downer
downier|downy
downiest|downy
dowy|dowie
dozier|dozy
doziest|dozy
drabber|drab
drabbest|drab
draftier|drafty
draftiest|drafty
draggier|draggy
draggiest|draggy
draughtier|draughty
draughtiest|draughty
dreamier|dreamy
dreamiest|dreamy
drearier|dreary
dreariest|dreary
dreggier|dreggy
dreggiest|dreggy
dresser|dresser
dressier|dressy
dressiest|dressy
drier|dry
driest|dry
drippier|drippy
drippiest|drippy
drowsier|drowsy
drowsiest|drowsy
dryer|dry
dryest|dry
dumpier|dumpy
dumpiest|dumpy
dunner|dun
dunnest|dun
duskier|dusky
duskiest|dusky
dustier|dusty
dustiest|dusty
earlier|early
earliest|early
earthier|earthy
earthiest|earthy
earthlier|earthly
earthliest|earthly
easier|easy
easiest|easy
easter|easter
eastsider|eastsider
edger|edger
edgier|edgy
edgiest|edgy
eerier|eerie
eeriest|eerie
emptier|empty
emptiest|empty
faker|faker
fancier|fancy
fanciest|fancy
fatter|fat
fattest|fat
fattier|fatty
fattiest|fatty
faultier|faulty
faultiest|faulty
feistier|feisty
feistiest|feisty
feller|feller
fiddlier|fiddly
fiddliest|fiddly
filmier|filmy
filmiest|filmy
filthier|filthy
filthiest|filthy
finnier|finny
finniest|finny
first-rater|first-rater
first-stringer|first-stringer
fishier|fishy
fishiest|fishy
fitter|fit
fittest|fit
flabbier|flabby
flabbiest|flabby
flaggier|flaggy
flaggiest|flaggy
flakier|flaky
flakiest|flaky
flasher|flasher
flashier|flashy
flashiest|flashy
flatter|flat
flattest|flat
flauntier|flaunty
flauntiest|flaunty
fledgier|fledgy
fledgiest|fledgy
fleecier|fleecy
fleeciest|fleecy
fleshier|fleshy
fleshiest|fleshy
fleshlier|fleshly
fleshliest|fleshly
flightier|flighty
flightiest|flighty
flimsier|flimsy
flimsiest|flimsy
flintier|flinty
flintiest|flinty
floatier|floaty
floatiest|floaty
floppier|floppy
floppiest|floppy
flossier|flossy
flossiest|flossy
fluffier|fluffy
fluffiest|fluffy
flukier|fluky
flukiest|fluky
foamier|foamy
foamiest|foamy
foggier|foggy
foggiest|foggy
folder|folder
folksier|folksy
folksiest|folksy
foolhardier|foolhardy
foolhardiest|foolhardy
fore-and-after|fore-and-after
foreigner|foreigner
forest|forest
founder|founder
foxier|foxy
foxiest|foxy
fratchier|fratchy
fratchiest|fratchy
freakier|freaky
freakiest|freaky
freer|free
freest|free
frenchier|frenchy
frenchiest|frenchy
friendlier|friendly
friendliest|friendly
friskier|frisky
friskiest|frisky
frizzier|frizzy
frizziest|frizzy
frizzlier|frizzly
frizzliest|frizzly
frostier|frosty
frostiest|frosty
frouzier|frouzy
frouziest|frouzy
frowsier|frowsy
frowsiest|frowsy
frowzier|frowzy
frowziest|frowzy
fruitier|fruity
fruitiest|fruity
funkier|funky
funkiest|funky
funnier|funny
funniest|funny
furrier|furry
furriest|furry
fussier|fussy
fussiest|fussy
fustier|fusty
fustiest|fusty
fuzzier|fuzzy
fuzziest|fuzzy
gabbier|gabby
gabbiest|gabby
gamier|gamy
gamiest|gamy
gammier|gammy
gammiest|gammy
gassier|gassy
gassiest|gassy
gaudier|gaudy
gaudiest|gaudy
gauzier|gauzy
gauziest|gauzy
gawkier|gawky
gawkiest|gawky
ghastlier|ghastly
ghastliest|ghastly
ghostlier|ghostly
ghostliest|ghostly
giddier|giddy
giddiest|giddy
gladder|glad
gladdest|glad
glassier|glassy
glassiest|glassy
glibber|glib
glibbest|glib
gloomier|gloomy
gloomiest|gloomy
glossier|glossy
glossiest|glossy
glummer|glum
glummest|glum
godlier|godly
godliest|godly
goer|goer
goner|goner
goodlier|goodly
goodliest|goodly
goofier|goofy
goofiest|goofy
gooier|gooey
gooiest|gooey
goosier|goosy
goosiest|goosy
gorier|gory
goriest|gory
gradelier|gradely
gradeliest|gradely
grader|grader
grainier|grainy
grainiest|grainy
grassier|grassy
grassiest|grassy
greasier|greasy
greasiest|greasy
greedier|greedy
greediest|greedy
grimmer|grim
grimmest|grim
grislier|grisly
grisliest|grisly
grittier|gritty
grittiest|gritty
grizzlier|grizzly
grizzliest|grizzly
groggier|groggy
groggiest|groggy
groovier|groovy
grooviest|groovy
grottier|grotty
grottiest|grotty
grounder|grounder
grouper|grouper
groutier|grouty
groutiest|grouty
grubbier|grubby
grubbiest|grubby
grumpier|grumpy
grumpiest|grumpy
guest|guest
guiltier|guilty
guiltiest|guilty
gummier|gummy
gummiest|gummy
gushier|gushy
gushiest|gushy
gustier|gusty
gustiest|gusty
gutsier|gutsy
gutsiest|gutsy
hairier|hairy
hairiest|hairy
halfways|halfway
halter|halter
hammier|hammy
hammiest|hammy
handier|handy
handiest|handy
happier|happy
happiest|happy
hardier|hardy
hardiest|hardy
hastier|hasty
hastiest|hasty
haughtier|haughty
haughtiest|haughty
hazier|hazy
haziest|hazy
header|header
headier|heady
headiest|heady
healthier|healthy
healthiest|healthy
heartier|hearty
heartiest|hearty
heavier|heavy
heaviest|heavy
heftier|hefty
heftiest|hefty
hepper|hep
heppest|hep
herbier|herby
herbiest|herby
hinder|hind
hipper|hip
hippest|hip
hippier|hippy
hippiest|hippy
hoarier|hoary
hoariest|hoary
holier|holy
holiest|holy
homelier|homely
homeliest|homely
homer|homer
homier|homey
homiest|homey
hornier|horny
horniest|horny
horsier|horsy
horsiest|horsy
hotter|hot
hottest|hot
humpier|humpy
humpiest|humpy
hunger|hunger
hungrier|hungry
hungriest|hungry
huskier|husky
huskiest|husky
icier|icy
iciest|icy
inkier|inky
inkiest|inky
insider|insider
interest|interest
jaggier|jaggy
jaggiest|jaggy
jammier|jammy
jammiest|jammy
jauntier|jaunty
jauntiest|jaunty
jazzier|jazzy
jazziest|jazzy
jerkier|jerky
jerkiest|jerky
jointer|jointer
jollier|jolly
jolliest|jolly
juicier|juicy
juiciest|juicy
jumpier|jumpy
jumpiest|jumpy
kindlier|kindly
kindliest|kindly
kinkier|kinky
kinkiest|kinky
knottier|knotty
knottiest|knotty
knurlier|knurly
knurliest|knurly
kookier|kooky
kookiest|kooky
lacier|lacy
laciest|lacy
lairier|lairy
lairiest|lairy
lakier|laky
lakiest|laky
lander|lander
lankier|lanky
lankiest|lanky
lathier|lathy
lathiest|lathy
layer|layer
lazier|lazy
laziest|lazy
leafier|leafy
leafiest|leafy
leakier|leaky
leakiest|leaky
learier|leary
leariest|leary
leerier|leery
leeriest|leery
leer|leer
left-hander|left-hander
left-winger|left-winger
leggier|leggy
leggiest|leggy
lengthier|lengthy
lengthiest|lengthy
ler|ler
leveler|leveler
limier|limy
limiest|limy
lippier|lippy
lippiest|lippy
liter|liter
livelier|lively
liveliest|lively
liver|liver
loather|loather
loftier|lofty
loftiest|lofty
logier|logy
logiest|logy
lonelier|lonely
loneliest|lonely
loner|loner
loonier|loony
looniest|loony
loopier|loopy
loopiest|loopy
lordlier|lordly
lordliest|lordly
lousier|lousy
lousiest|lousy
lovelier|lovely
loveliest|lovely
lowlander|lowlander
lowlier|lowly
lowliest|lowly
luckier|lucky
luckiest|lucky
lumpier|lumpy
lumpiest|lumpy
lunier|luny
luniest|luny
lustier|lusty
lustiest|lusty
madder|mad
maddest|mad
mainer|mainer
maligner|maligner
maltier|malty
maltiest|malty
mangier|mangy
mangiest|mangy
mankier|manky
mankiest|manky
manlier|manly
manliest|manly
mariner|mariner
marshier|marshy
marshiest|marshy
massier|massy
massiest|massy
matter|matter
maungier|maungy
maungiest|maungy
mazier|mazy
maziest|mazy
mealier|mealy
mealiest|mealy
measlier|measly
measliest|measly
meatier|meaty
meatiest|meaty
meeter|meeter
merrier|merry
merriest|merry
messier|messy
messiest|messy
miffier|miffy
miffiest|miffy
mightier|mighty
mightiest|mighty
milcher|milcher
milker|milker
milkier|milky
milkiest|milky
mingier|mingy
mingiest|mingy
minter|minter
mirkier|mirky
mirkiest|mirky
miser|miser
mistier|misty
mistiest|misty
mocker|mocker
modeler|modeler
modest|modest
moldier|moldy
moldiest|moldy
moodier|moody
moodiest|moody
moonier|moony
mooniest|moony
mothier|mothy
mothiest|mothy
mouldier|mouldy
mouldiest|mouldy
mousier|mousy
mousiest|mousy
mouthier|mouthy
mouthiest|mouthy
muckier|mucky
muckiest|mucky
muddier|muddy
muddiest|muddy
muggier|muggy
muggiest|muggy
multiplexer|multiplexer
murkier|murky
murkiest|murky
mushier|mushy
mushiest|mushy
muskier|musky
muskiest|musky
muster|muster
mustier|musty
mustiest|musty
muzzier|muzzy
muzziest|muzzy
nappier|nappy
nappiest|nappy
nastier|nasty
nastiest|nasty
nattier|natty
nattiest|natty
naughtier|naughty
naughtiest|naughty
needier|needy
neediest|needy
nervier|nervy
nerviest|nervy
newsier|newsy
newsiest|newsy
niftier|nifty
niftiest|nifty
nippier|nippy
nippiest|nippy
nittier|nitty
nittiest|nitty
noisier|noisy
noisiest|noisy
northeasterner|northeasterner
northerner|northerner
norther|norther
nosier|nosy
nosiest|nosy
number|number
nuttier|nutty
nuttiest|nutty
offer|offer
oilier|oily
oiliest|oily
old-timer|old-timer
oliver|oliver
oozier|oozy
ooziest|oozy
opener|opener
outsider|outsider
overcomer|overcomer
overnighter|overnighter
owner|owner
pallier|pally
palliest|pally
palmier|palmy
palmiest|palmy
paltrier|paltry
paltriest|paltry
pappier|pappy
pappiest|pappy
parkier|parky
parkiest|parky
part-timer|part-timer
passer|passer
paster|paster
pastier|pasty
pastiest|pasty
patchier|patchy
patchiest|patchy
pater|pater
pawkier|pawky
pawkiest|pawky
peachier|peachy
peachiest|peachy
pearler|pearler
pearlier|pearly
pearliest|pearly
pedaler|pedaler
peppier|peppy
peppiest|peppy
perkier|perky
perkiest|perky
peskier|pesky
peskiest|pesky
peter|peter
pettier|petty
pettiest|petty
phonier|phony
phoniest|phony
pickier|picky
pickiest|picky
piggier|piggy
piggiest|piggy
pinier|piny
piniest|piny
pitchier|pitchy
pitchiest|pitchy
pithier|pithy
pithiest|pithy
planer|planer
plashier|plashy
plashiest|plashy
platier|platy
platiest|platy
player|player
pluckier|plucky
pluckiest|plucky
plumber|plumber
plumier|plumy
plumiest|plumy
plummier|plummy
plummiest|plummy
podgier|podgy
podgiest|podgy
pokier|poky
pokiest|poky
polisher|polisher
porkier|porky
porkiest|porky
porter|porter
portlier|portly
portliest|portly
poster|poster
pottier|potty
pottiest|potty
preachier|preachy
preachiest|preachy
presenter|presenter
pretender|pretender
prettier|pretty
prettiest|pretty
pricier|pricy
priciest|pricy
pricklier|prickly
prickliest|prickly
priestlier|priestly
priestliest|priestly
primer|primer
primmer|prim
primmest|prim
princelier|princely
princeliest|princely
printer|printer
prissier|prissy
prissiest|prissy
privateer|privateer
privier|privy
priviest|privy
prompter|prompter
prosier|prosy
prosiest|prosy
pudgier|pudgy
pudgiest|pudgy
puffer|puffer
puffier|puffy
puffiest|puffy
pulpier|pulpy
pulpiest|pulpy
punchier|punchy
punchiest|punchy
punier|puny
puniest|puny
pushier|pushy
pushiest|pushy
pussier|pussy
pussiest|pussy
quaggier|quaggy
quaggiest|quaggy
quakier|quaky
quakiest|quaky
queasier|queasy
queasiest|queasy
queenlier|queenly
queenliest|queenly
racier|racy
raciest|racy
rainier|rainy
rainiest|rainy
randier|randy
randiest|randy
rangier|rangy
rangiest|rangy
ranker|ranker
rattier|ratty
rattiest|ratty
rattlier|rattly
rattliest|rattly
raunchier|raunchy
raunchiest|raunchy
readier|ready
readiest|ready
recorder|recorder
redder|red
reddest|red
reedier|reedy
reediest|reedy
renter|renter
retailer|retailer
right-hander|right-hander
right-winger|right-winger
rimier|rimy
rimiest|rimy
riskier|risky
riskiest|risky
ritzier|ritzy
ritziest|ritzy
roaster|roaster
rockier|rocky
rockiest|rocky
roilier|roily
roiliest|roily
rookier|rooky
rookiest|rooky
roomier|roomy
roomiest|roomy
ropier|ropy
ropiest|ropy
rosier|rosy
rosiest|rosy
rowdier|rowdy
rowdiest|rowdy
ruddier|ruddy
ruddiest|ruddy
runnier|runny
runniest|runny
rusher|rusher
rushier|rushy
rushiest|rushy
rustier|rusty
rustiest|rusty
ruttier|rutty
ruttiest|rutty
sadder|sad
saddest|sad
salter|salter
saltier|salty
saltiest|salty
sampler|sampler
sandier|sandy
sandiest|sandy
sappier|sappy
sappiest|sappy
sassier|sassy
sassiest|sassy
saucier|saucy
sauciest|saucy
savvier|savvy
savviest|savvy
scabbier|scabby
scabbiest|scabby
scalier|scaly
scaliest|scaly
scantier|scanty
scantiest|scanty
scarier|scary
scariest|scary
scraggier|scraggy
scraggiest|scraggy
scragglier|scraggly
scraggliest|scraggly
scraper|scraper
scrappier|scrappy
scrappiest|scrappy
scrawnier|scrawny
scrawniest|scrawny
screwier|screwy
screwiest|screwy
scrubbier|scrubby
scrubbiest|scrubby
scruffier|scruffy
scruffiest|scruffy
scungier|scungy
scungiest|scungy
scurvier|scurvy
scurviest|scurvy
seamier|seamy
seamiest|seamy
second-rater|second-rater
seconder|seconder
seedier|seedy
seediest|seedy
seemlier|seemly
seemliest|seemly
serer|serer
sexier|sexy
sexiest|sexy
shabbier|shabby
shabbiest|shabby
shadier|shady
shadiest|shady
shaggier|shaggy
shaggiest|shaggy
shakier|shaky
shakiest|shaky
shapelier|shapely
shapeliest|shapely
shier|shy
shiest|shy
shiftier|shifty
shiftiest|shifty
shinier|shiny
shiniest|shiny
shirtier|shirty
shirtiest|shirty
shoddier|shoddy
shoddiest|shoddy
showier|showy
showiest|showy
shrubbier|shrubby
shrubbiest|shrubby
shyer|shy
shyest|shy
sicklier|sickly
sickliest|sickly
sightlier|sightly
sightliest|sightly
signaler|signaler
signer|signer
silkier|silky
silkiest|silky
sillier|silly
silliest|silly
sketchier|sketchy
sketchiest|sketchy
skewer|skewer
skimpier|skimpy
skimpiest|skimpy
skinnier|skinny
skinniest|skinny
slaphappier|slaphappy
slaphappiest|slaphappy
slatier|slaty
slatiest|slaty
slaver|slaver
sleazier|sleazy
sleaziest|sleazy
sleepier|sleepy
sleepiest|sleepy
slier|sly
sliest|sly
slimier|slimy
slimiest|slimy
slimmer|slim
slimmest|slim
slimsier|slimsy
slimsiest|slimsy
slinkier|slinky
slinkiest|slinky
slippier|slippy
slippiest|slippy
sloppier|sloppy
sloppiest|sloppy
slyer|sly
slyest|sly
smarmier|smarmy
smarmiest|smarmy
smellier|smelly
smelliest|smelly
smokier|smoky
smokiest|smoky
smugger|smug
smuggest|smug
snakier|snaky
snakiest|snaky
snappier|snappy
snappiest|snappy
snatchier|snatchy
snatchiest|snatchy
snazzier|snazzy
snazziest|snazzy
sneaker|sneaker
sniffier|sniffy
sniffiest|sniffy
snootier|snooty
snootiest|snooty
snottier|snotty
snottiest|snotty
snowier|snowy
snowiest|snowy
snuffer|snuffer
snuffier|snuffy
snuffiest|snuffy
snugger|snug
snuggest|snug
soapier|soapy
soapiest|soapy
soggier|soggy
soggiest|soggy
solder|solder
sonsier|sonsy
sonsiest|sonsy
sootier|sooty
sootiest|sooty
soppier|soppy
soppiest|soppy
sorrier|sorry
sorriest|sorry
soupier|soupy
soupiest|soupy
southerner|southerner
souther|souther
speedier|speedy
speediest|speedy
spicier|spicy
spiciest|spicy
spiffier|spiffy
spiffiest|spiffy
spikier|spiky
spikiest|spiky
spindlier|spindly
spindliest|spindly
spinier|spiny
spiniest|spiny
splashier|splashy
splashiest|splashy
spongier|spongy
spongiest|spongy
spookier|spooky
spookiest|spooky
spoonier|spoony
spooniest|spoony
sportier|sporty
sportiest|sporty
spottier|spotty
spottiest|spotty
spreader|spreader
sprier|spry
spriest|spry
sprightlier|sprightly
sprightliest|sprightly
springer|springer
springier|springy
springiest|springy
squashier|squashy
squashiest|squashy
squatter|squat
squattest|squat
squattier|squatty
squattiest|squatty
squiffier|squiffy
squiffiest|squiffy
stagier|stagy
stagiest|stagy
stalkier|stalky
stalkiest|stalky
stapler|stapler
starchier|starchy
starchiest|starchy
starer|starer
starest|starest
starrier|starry
starriest|starry
statelier|stately
stateliest|stately
steadier|steady
steadiest|steady
stealthier|stealthy
stealthiest|stealthy
steamier|steamy
steamiest|steamy
stingier|stingy
stingiest|stingy
stiper|striper
stocker|stocker
stockier|stocky
stockiest|stocky
stodgier|stodgy
stodgiest|stodgy
stonier|stony
stoniest|stony
stormier|stormy
stormiest|stormy
streakier|streaky
streakiest|streaky
streamier|streamy
streamiest|streamy
stretcher|stretcher
stretchier|stretchy
stretchiest|stretchy
stringier|stringy
stringiest|stringy
stripier|stripy
stripiest|stripy
stronger|strong
strongest|strong
stroppier|stroppy
stroppiest|stroppy
stuffier|stuffy
stuffiest|stuffy
stumpier|stumpy
stumpiest|stumpy
sturdier|sturdy
sturdiest|sturdy
submariner|submariner
sulkier|sulky
sulkiest|sulky
sultrier|sultry
sultriest|sultry
sunnier|sunny
sunniest|sunny
surlier|surly
surliest|surly
swagger|swagger
swankier|swanky
swankiest|swanky
swarthier|swarthy
swarthiest|swarthy
sweatier|sweaty
sweatiest|sweaty
tackier|tacky
tackiest|tacky
talkier|talky
talkiest|talky
tangier|tangy
tangiest|tangy
tanner|tan
tannest|tan
tardier|tardy
tardiest|tardy
tastier|tasty
tastiest|tasty
tattier|tatty
tattiest|tatty
tawdrier|tawdry
tawdriest|tawdry
techier|techy
techiest|techy
teenager|teenager
teenier|teeny
teeniest|teeny
teetotaler|teetotaler
tester|tester
testier|testy
testiest|testy
tetchier|tetchy
tetchiest|tetchy
thinner|thin
thinnest|thin
third-rater|third-rater
thirstier|thirsty
thirstiest|thirsty
thornier|thorny
thorniest|thorny
threadier|thready
threadiest|thready
thriftier|thrifty
thriftiest|thrifty
throatier|throaty
throatiest|throaty
tidier|tidy
tidiest|tidy
timelier|timely
timeliest|timely
tinier|tiny
tiniest|tiny
tinnier|tinny
tinniest|tinny
tipsier|tipsy
tipsiest|tipsy
tonier|tony
toniest|tony
toothier|toothy
toothiest|toothy
toper|toper
touchier|touchy
touchiest|touchy
trader|trader
trashier|trashy
trashiest|trashy
trendier|trendy
trendiest|trendy
trickier|tricky
trickiest|tricky
tricksier|tricksy
tricksiest|tricksy
trimer|trimer
trimmer|trim
trimmest|trim
truer|true
truest|true
trustier|trusty
trustiest|trusty
tubbier|tubby
tubbiest|tubby
turfier|turfy
turfiest|turfy
tweedier|tweedy
tweediest|tweedy
twiggier|twiggy
twiggiest|twiggy
uglier|ugly
ugliest|ugly
unfriendlier|unfriendly
unfriendliest|unfriendly
ungainlier|ungainly
ungainliest|ungainly
ungodlier|ungodly
ungodliest|ungodly
unhappier|unhappy
unhappiest|unhappy
unhealthier|unhealthy
unhealthiest|unhealthy
unholier|unholy
unholiest|unholy
unrulier|unruly
unruliest|unruly
untidier|untidy
untidiest|untidy
vastier|vasty
vastiest|vasty
vest|vest
viewier|viewy
viewiest|viewy
wackier|wacky
wackiest|wacky
wanner|wan
wannest|wan
warier|wary
wariest|wary
washier|washy
washiest|washy
waster|waster
wavier|wavy
waviest|wavy
waxier|waxy
waxiest|waxy
weaklier|weakly
weakliest|weakly
wealthier|wealthy
wealthiest|wealthy
wearier|weary
weariest|weary
webbier|webby
webbiest|webby
weedier|weedy
weediest|weedy
weenier|weeny
weeniest|weeny
weensier|weensy
weensiest|weensy
weepier|weepy
weepiest|weepy
weightier|weighty
weightiest|weighty
well|good
welsher|welsher
wetter|wet
wettest|wet
whackier|whacky
whackiest|whacky
whimsier|whimsy
whimsiest|whimsy
wholesaler|wholesaler
wieldier|wieldy
wieldiest|wieldy
wilier|wily
wiliest|wily
windier|windy
windiest|windy
winier|winy
winiest|winy
winterier|wintery
winteriest|wintery
wintrier|wintry
wintriest|wintry
wirier|wiry
wiriest|wiry
wispier|wispy
wispiest|wispy
wittier|witty
wittiest|witty
wonkier|wonky
wonkiest|wonky
woodier|woody
woodiest|woody
woodsier|woodsy
woodsiest|woodsy
woollier|woolly
woolliest|woolly
woozier|woozy
wooziest|woozy
wordier|wordy
wordiest|wordy
worldlier|worldly
worldliest|worldly
wormier|wormy
wormiest|wormy
worse|bad
worst|bad
worthier|worthy
worthiest|worthy
wrier|wry
wriest|wry
wryer|wry
wryest|wry
yarer|yare
yarest|yare
yeastier|yeasty
yeastiest|yeasty
younger|young
youngest|young
yummier|yummy
yummiest|yummy
zanier|zany
zaniest|zany
zippier|zippy
zippiest|zippy