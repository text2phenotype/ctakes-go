er|
est|
er|e
est|e