'd|have
'mmm|be
'm|be
're|be
've|have
abetted|abet
abetting|abet
abhorred|abhor
abhorring|abhor
abode|abide
abought|aby
about-shipped|about-ship
about-shipping|about-ship
abutted|abut
abutting|abut
abye|aby
accompanied|accompany
acetified|acetify
acidified|acidify
acquitted|acquit
acquitting|acquit
ad-libbed|ad-lib
ad-libbing|ad-lib
addrest|address
admitted|admit
admitting|admit
aerified|aerify
air-dried|air-dry
airdropped|airdrop
airdropping|airdrop
alkalified|alkalify
allied|ally
allotted|allot
allotting|allot
allowed_for|allow_for
allowing_for|allow_for
allows_for|allow_for
ammonified|ammonify
amnestied|amnesty
amplified|amplify
am|be
anglified|anglify
annulled|annul
annulling|annul
appalled|appal
appalling|appal
appall|appal
applied|apply
arcked|arc
arcking|arc
are|be
argufied|argufy
arisen|arise
arose|arise
ate|eat
atrophied|atrophy
averred|aver
averring|aver
awoken|awake
awoke|awake
babied|baby
baby-sat|baby-sit
baby-sitting|baby-sit
back-pedalled|back-pedal
back-pedalling|back-pedal
backbitten|backbite
backbit|backbite
backslidden|backslide
backslid|backslide
bade|bid
bagged|bag
bagging|bag
ballyragged|ballyrag
ballyragging|ballyrag
bandied|bandy
banned|ban
banning|ban
barred|bar
barrelled|barrel
barrelling|barrel
barring|bar
basified|basify
batted|bat
batting|bat
bayonetted|bayonet
bayonetting|bayonet
beaten|beat
beatified|beatify
beautified|beautify
became_known|become_known
became|become
becomes_known|become_known
bedded|bed
bedding|bed
bedevilled|bedevil
bedevilling|bedevil
bedimmed|bedim
bedimming|bedim
bed|bed
been|be
befallen|befall
befell|befall
befitted|befit
befitting|befit
befogged|befog
befogging|befog
began|begin
begat|beget
begetting|beget
begged|beg
begging|beg
beginning|begin
begirt|begird
begotten|beget
begot|beget
begun|begin
beheld|behold
beholden|behold
bejewelled|bejewel
bejewelling|bejewel
bellied|belly
belly-flopped|belly-flop
belly-flopping|belly-flop
belying|belie
benefitted|benefit
benefitting|benefit
benempt|bename
bent|bend
berried|berry
besetting|beset
besought|beseech
bespoken|bespeak
bespoke|bespeak
bestirred|bestir
bestirring|bestir
bestrewn|bestrew
bestridden|bestride
bestrid|bestride
bestrode|bestride
betaken|betake
bethought|bethink
betook|betake
betted|bet
betting|bet
bevelled|bevel
bevelling|bevel
biassed|bias
biassing|bias
bidden|bid
bidding|bid
bing|bing
binned|bin
binning|bin
bird-dogged|bird-dog
bird-dogging|bird-dog
bitted|bit
bitten|bite
bitting|bit
bit|bite
bivouacked|bivouac
bivouacking|bivouac
blabbed|blab
blabbing|blab
blackberried|blackberry
blacklegged|blackleg
blacklegging|blackleg
blatted|blat
blatting|blat
bled|bleed
blest|bless
blew_one's_nose|blow_one's_nose
blew|blow
blipped|blip
blipping|blip
blobbed|blob
blobbing|blob
bloodied|bloody
blotted|blot
blotting|blot
blowing_one's_nose|blow_one's_nose
blown|blow
blows_one's_nose|blow_one's_nose
blubbed|blub
blubbing|blub
blue-pencilled|blue-pencil
blue-pencilling|blue-pencil
blurred|blur
blurring|blur
bobbed|bob
bobbing|bob
bodied|body
bogged-down|bog-down
bogged_down|bog_down
bogged|bog
bogging-down|bog-down
bogging_down|bog_down
bogging|bog
bogs-down|bog-down
bogs_down|bog_down
bondin'|bond
booby-trapped|booby-trap
booby-trapping|booby-trap
bootlegged|bootleg
bootlegging|bootleg
bopped|bop
bopping|bop
bore|bear
borne|bear
born|bear
bottle-fed|bottle-feed
bought|buy
bound|bind
bragged|brag
bragging|brag
breast-fed|breast-feed
bred|breed
brevetted|brevet
brevetting|brevet
brimmed|brim
brimming|brim
broken|break
broke|break
brought|bring
browbeaten|browbeat
brutified|brutify
budded|bud
budding|bud
bugged|bug
bugging|bug
built|build
bulldogging|bulldog
bullied|bully
bullshitted|bullshit
bullshitting|bullshit
bullwhipped|bullwhip
bullwhipping|bullwhip
bullyragged|bullyrag
bullyragging|bullyrag
bummed|bum
bumming|bum
buried|bury
burnt|burn
burred|bur
burring|bur
bushelled|bushel
bushelling|bushel
busied|busy
bypast|bypass
caballed|cabal
caballing|cabal
caddied|caddie
caddies|caddie
caddying|caddie
caddy|caddie
calcified|calcify
came|come
canalled|canal
canalling|canal
cancelled|cancel
cancelling|cancel
candied|candy
canned|can
canning|can
canopied|canopy
capped|cap
capping|cap
carburetted|carburet
carburetting|carburet
carillonned|carillon
carillonning|carillon
carnied|carny
carnified|carnify
carolled|carol
carolling|carol
carried|carry
casefied|casefy
catnapped|catnap
catnapping|catnap
catted|cat
catting|cat
caught|catch
cavilled|cavil
cavilling|cavil
certified|certify
channelled|channel
channelling|channel
chapped|chap
chapping|chap
charred|char
charring|char
chatted|chat
chatting|chat
chevied|chivy
chevies|chivy
chevying|chivy
chidden|chide
chid|chide
chinned|chin
chinning|chin
chipped|chip
chipping|chip
chiselled|chisel
chiselling|chisel
chitchatted|chitchat
chitchatting|chitchat
chivied|chivy
chivved|chiv
chivvied|chivy
chivvies|chivy
chivving|chiv
chivvying|chivy
chondrified|chondrify
chopped|chop
chopping|chop
chosen|choose
chose|choose
chugged|chug
chugging|chug
chummed|chum
chumming|chum
citified|citify
cladding|clad
clad|clothe
clammed|clam
clamming|clam
clapped|clap
clapping|clap
clarified|clarify
classified|classify
cleft|cleave
clemmed|clem
clemming|clem
clept|clepe
clipped|clip
clipping|clip
clogged|clog
clogging|clog
clopped|clop
clopping|clop
clotted|clot
clotting|clot
cloven|cleave
clove|cleave
clubbed|club
clubbing|club
clung|cling
co-opted|coopt
co-opting|coopt
co-opts|coopts
co-ordinated|coordinate
co-ordinates|coordinate
co-ordinate|coordinate
co-ordinating|coordinate
co-starred|co-star
co-starring|co-star
cockneyfied|cockneyfy
codded|cod
codding|cod
codified|codify
cogged|cog
cogging|cog
coiffed|coif
coiffing|coif
collied|colly
combatted|combat
combatting|combat
committed|commit
committing|commit
compelled|compel
compelling|compel
complied|comply
complotted|complot
complotting|complot
concurred|concur
concurring|concur
confabbed|confab
confabbing|confab
conferred|confer
conferring|confer
conned|con
conning|con
controlled|control
controlling|control
copied|copy
copped|cop
copping|cop
coquetted|coquet
coquetting|coquet
corralled|corral
corralling|corral
counselled|counsel
counselling|counsel
counterplotted|counterplot
counterplotting|counterplot
countersank|countersink
countersunk|countersink
court-martialled|court-martial
court-martialling|court-martial
coverred|cover
crabbed|crab
crabbing|crab
crammed|cram
cramming|cram
crapped|crap
crapping|crap
crept|creep
cribbed|crib
cribbing|crib
cried|cry
cropped|crop
cropping|crop
crossbred|crossbreed
crosscutting|crosscut
crucified|crucify
cubbed|cub
cubbing|cub
cudgelled|cudgel
cudgelling|cudgel
cupelled|cupel
cupelling|cupel
cupped|cup
cupping|cup
curetted|curet
curettes|curet
curetting|curet
curried|curry
curst|curse
curtsied|curtsy
curvetted|curvet
curvetting|curvet
cutting|cut
dabbed|dab
dabbing|dab
dagged|dag
dagging|dag
dallied|dally
dammed|dam
damming|dam
damnified|damnify
dandified|dandify
dapped|dap
dapping|dap
dealt|deal
debarred|debar
debarring|debar
debugged|debug
debugging|debug
debussed|debus
debusses|debus
debussing|debus
decalcified|decalcify
declassified|declassify
decontrolled|decontrol
decontrolling|decontrol
decried|decry
deep-freezed|deepfreeze
deep-freezes|deepfreeze
deep-freeze|deepfreeze
deep-fried|deep-fry
deferred|defer
deferring|defer
defied|defy
degassed|degas
degasses|degas
degassing|degas
dehumidified|dehumidify
deified|deify
demitted|demit
demitting|demit
demobbed|demob
demobbing|demob
demulsified|demulsify
demurred|demur
demurring|demur
demystified|demystify
denazified|denazify
denied|deny
denitrified|denitrify
denned|den
denning|den
descried|descry
deterred|deter
deterring|deter
detoxified|detoxify
devilled|devil
devilling|devil
devitrified|devitrify
diagrammed|diagram
diagramming|diagram
dialled|dial
dialling|dial
dibbed|dib
dibbing|dib
did|do
digging|dig
dignified|dignify
dilly-dallied|dilly-dally
dimmed|dim
dimming|dim
dinned|din
dinning|din
dipped|dip
dipping|dip
dirtied|dirty
disannulled|disannul
disannulling|disannul
disbarred|disbar
disbarring|disbar
disbudded|disbud
disbudding|disbud
disembodied|disembody
disembowelled|disembowel
disembowelling|disembowel
disenthralled|disenthral
disenthralling|disenthral
disenthralls|disenthral
disenthrall|disenthral
disenthrals|disenthrall
dishevelled|dishevel
dishevelling|dishevel
disinterred|disinter
disinterring|disinter
dispelled|dispel
dispelling|dispel
disproven|disprove
disqualified|disqualify
dissatisfied|dissatisfy
distilled|distil
distilling|distil
distill|distil
diversified|diversify
divvied|divvy
dizzied|dizzy
dogged|dog
dogging|dog
doglegged|dogleg
doglegging|dogleg
dollied|dolly
done|do
donned|don
donning|don
dotted|dot
dotting|dot
dought|dow
dove|dive
drabbed|drab
drabbing|drab
dragged|drag
dragging|drag
drank|drink
drawn|draw
dreamt|dream
drew|draw
dried|dry
dripped|drip
dripping|drip
drivelled|drivel
drivelling|drivel
driven|drive
dropped|drop
dropping|drop
drove|drive
drubbed|drub
drubbing|drub
drugged|drug
drugging|drug
drummed|drum
drumming|drum
drunk|drink
dubbed|dub
dubbing|dub
duelled|duel
duelling|duel
dug|dig
dulcified|dulcify
dummied|dummy
dunned|dun
dunning|dun
dwelt|dwell
dying|die
e-mailed|email
e-mailing|email
e-mail|email
easied|easy
eaten|eat
eavesdropped|eavesdrop
eavesdropping|eavesdrop
eddied|eddy
edified|edify
ego-tripped|ego-trip
ego-tripping|ego-trip
electrified|electrify
embedded|embed
embedding|embed
embodied|embody
embussed|embus
embusses|embus
embussing|embus
emitted|emit
emitting|emit
empanelled|empanel
empanelling|empanel
emptied|empty
emulsified|emulsify
enamelled|enamel
enamelling|enamel
englutted|englut
englutting|englut
enrolled|enrol
enrolling|enrol
enroll|enrol
enthralled|enthral
enthralling|enthral
enthrall|enthral
entrammelled|entrammel
entrammelling|entrammel
entrapped|entrap
entrapping|entrap
envied|envy
enwound|enwind
enwrapped|enwrap
enwrapping|enwrap
equalled|equal
equalling|equal
equipped|equip
equipping|equip
espied|espy
esterified|esterify
estopped|estop
estopping|estop
etherified|etherify
excelled|excel
excelling|excel
exemplified|exemplify
expelled|expel
expelling|expel
extolled|extol
extolling|extol
extoll|extol
facetted|facet
facetting|facet
fagged|fag
fagging|fag
fallen|fall
falsified|falsify
fancied|fancy
fanned|fan
fanning|fan
fantasied|fantasy
fatted|fat
fatting|fat
featherbedded|featherbed
featherbedding|featherbed
fed|feed
feed|feed
fee|feed
fell|fall
felt|feel
ferried|ferry
fibbed|fib
fibbing|fib
figged|fig
figging|fig
filled_up|fill_up
fine-drawn|fine-draw
fine-drew|fine-draw
finned|fin
finning|fin
fitted|fit
fitting|fit
flagged|flag
flagging|flag
flammed|flam
flamming|flam
flannelled|flannel
flannelling|flannel
flapped|flap
flapping|flap
flatted|flat
flatting|flat
fled|flee
flew|fly
flimflammed|flimflam
flimflamming|flimflam
flip-flopped|flip-flop
flip-flopping|flip-flop
flipped|flip
flipping|flip
flitted|flit
flitting|flit
flogged|flog
flogging|flog
floodlit|floodlight
flopped|flop
flopping|flop
flown|fly
flubbed|flub
flubbing|flub
flung|fling
flurried|flurry
flyblew|flyblow
flyblown|flyblow
fobbed|fob
fobbing|fob
focussed|focus
fogged|fog
fogging|fog
footslogged|footslog
footslogging|footslog
forbade|forbid
forbad|forbid
forbidden|forbid
forbidding|forbid
forbore|forbear
forborne|forbear
force-fed|force-feed
fordid|fordo
fordone|fordo
foredid|foredo
foredone|foredo
foregone|forego
foreknew|foreknow
foreknown|foreknow
foreran|forerun
forerunning|forerun
foresaw|foresee
foreseen|foresee
foreshown|foreshow
forespoken|forespeak
forespoke|forespeak
foretold|foretell
forewent|forego
forgave|forgive
forgetting|forget
forgiven|forgive
forgone|forgo
forgotten|forget
forgot|forget
formatted|format
formatting|format
forsaken|forsake
forsook|forsake
forspoken|forspeak
forspoke|forspeak
forswore|forswear
forsworn|forswear
fortified|fortify
forwent|forgo
fought|fight
found|find
foxtrotted|foxtrot
foxtrotting|foxtrot
frapped|frap
frapping|frap
freeze-dried|freeze-dry
frenchified|frenchify
frenzied|frenzy
fretted|fret
fretting|fret
fried|fry
frigged|frig
frigging|frig
fritted|frit
fritting|frit
fritt|frit
frivolled|frivol
frivolling|frivol
frogged|frog
frogging|frog
frolicked|frolic
frolicking|frolic
frozen|freeze
froze|freeze
fructified|fructify
fuelled|fuel
fuelling|fuel
fulfilled|fulfil
fulfilling|fulfil
fulfill|fulfil
funned|fun
funnelled|funnel
funnelling|funnel
funning|fun
furred|fur
furring|fur
gadded|gad
gadding|gad
gagged|gag
gagging|gag
gainsaid|gainsay
gambolled|gambol
gambolling|gambol
gammed|gam
gamming|gam
ganned|gan
ganning|gan
gan|gin
gapped|gap
gapping|gap
gasified|gasify
gassed|gas
gasses|gas
gassing|gas
gave|give
gelled|gel
gelling|gel
gelt|geld
gemmed|gem
gemming|gem
genned-up|gen-up
genning-up|gen-up
gens-up|gen-up
gets_lost|get_lost
gets_started|get_started
getting_lost|get_lost
getting_started|get_started
getting|get
ghostwritten|ghostwrite
ghostwrote|ghostwrite
gibbed|gib
gibbing|gib
giddied|giddy
giftwrapped|giftwrap
giftwrapping|giftwrap
gigged|gig
gigging|gig
gilt|gild
ginned|gin
ginning|gin
gipped|gip
gipping|gip
girt|gird
given|give
glommed|glom
glomming|glom
gloried|glory
glorified|glorify
glutted|glut
glutting|glut
gnawn|gnaw
goes_deep|go_deep
going_deep|go_deep
gollied|golly
gone_deep|go_deep
gone|go
goose-stepped|goose-step
goose-stepping|goose-step
got_lost|get_lost
got_started|get_started
gotten_lost|get_lost
gotten|get
got|get
grabbed|grab
grabbing|grab
gratified|gratify
gravelled|gravel
gravelling|gravel
graven|grave
grew|grow
grinned|grin
grinning|grin
gripped|grip
gripping|grip
gript|grip
gritted|grit
gritting|grit
ground|grind
grovelled|grovel
grovelling|grovel
grown|grow
grubbed|grub
grubbing|grub
guarantied|guaranty
gullied|gully
gummed|gum
gumming|gum
gunned|gun
gunning|gun
gypped|gyp
gypping|gyp
hacksawn|hacksaw
had_a_feeling|have_a_feeling
had_left|have_left
had_the_feeling|have_the_feeling
had|have
hammed|ham
hamming|ham
hamstrung|hamstring
hand-knitted|hand-knit
hand-knitting|hand-knit
handfed|handfeed
handicapped|handicap
handicapping|handicap
handselled|handsel
handselling|handsel
harried|harry
has_a_feeling|have_a_feeling
has_left|have_left
has_the_feeling|have_the_feeling
has|have
hatchelled|hatchel
hatchelling|hatchel
hatted|hat
hatting|hat
having_a_feeling|have_a_feeling
having_left|have_left
having_the_feeling|have_the_feeling
heard|hear
hedgehopped|hedgehop
hedgehopping|hedgehop
held|hold
hemmed|hem
hemming|hem
hewn|hew
hiccupped|hiccup
hiccupping|hiccup
hidden|hide
hid|hide
high-hatted|high-hat
high-hatting|high-hat
hinnied|hinny
hitting|hit
hobbed|hob
hobbing|hob
hobnobbed|hobnob
hobnobbing|hobnob
hocus-pocussed|hocus-pocus
hocus-pocussing|hocus-pocus
hocussed|hocus
hocussing|hocus
hogged|hog
hogging|hog
hogtying|hogtie
honied|honey
hopped|hop
hopping|hop
horrified|horrify
horsewhipped|horsewhip
horsewhipping|horsewhip
houselled|housel
houselling|housel
hovelled|hovel
hovelling|hovel
hove|heave
hugged|hug
hugging|hug
humbugged|humbug
humbugging|humbug
humidified|humidify
hummed|hum
humming|hum
hung|hang
hurried|hurry
hypertrophied|hypertrophy
identified|identify
imbedded|imbed
imbedding|imbed
impanelled|impanel
impanelling|impanel
impelled|impel
impelling|impel
implied|imply
inbred|inbreed
incurred|incur
incurring|incur
indemnified|indemnify
indwelt|indwell
inferred|infer
inferring|infer
initialled|initial
initialling|initial
inlaid|inlay
insetting|inset
inspanned|inspan
inspanning|inspan
installed|instal
installing|instal
install|instal
intensified|intensify
interbred|interbreed
intercropped|intercrop
intercropping|intercrop
intercutting|intercut
interlaid|interlay
interlapped|interlap
interlapping|interlap
intermarried|intermarry
intermitted|intermit
intermitting|intermit
interpled|interplead
interred|inter
interring|inter
interstratified|interstratify
interwoven|interweave
interwove|interweave
intromitted|intromit
intromitting|intromit
inwoven|inweave
inwove|inweave
inwrapped|inwrap
inwrapping|inwrap
is|be
jabbed|jab
jabbing|jab
jagged|jag
jagging|jag
jammed|jam
jamming|jam
japanned|japan
japanning|japan
jarred|jar
jarring|jar
jellied|jelly
jellified|jellify
jemmied|jemmy
jerry-built|jerry-build
jetted|jet
jetting|jet
jewelled|jewel
jewelling|jewel
jibbed|jib
jibbing|jib
jigged|jig
jigging|jig
jimmied|jimmy
jitterbugged|jitterbug
jitterbugging|jitterbug
jobbed|job
jobbing|job
jog-trotted|jog-trot
jog-trotting|jog-trot
jogged|jog
jogging|jog
joined_battle|join_battle
joined_forces|join_forces
joining_battle|join_battle
joining_forces|join_forces
joins_battle|join_battle
joins_forces|join_forces
jollied|jolly
jollified|jollify
jotted|jot
jotting|jot
joy-ridden|joy-ride
joy-rode|joy-ride
joypopped|joypop
joypopping|joypop
jugged|jug
jugging|jug
jumped_off|jump_off
jumping_off|jump_off
jumps_off|jump_off
justified|justify
jutted|jut
jutting|jut
kenned|ken
kennelled|kennel
kennelling|kennel
kenning|ken
kent|ken
kept|keep
kernelled|kernel
kernelling|kernel
kidded|kid
kidding|kid
kidnapped|kidnap
kidnapping|kidnap
kipped|kip
kipping|kip
knapped|knap
knapping|knap
kneecapped|kneecap
kneecapping|kneecap
knelt|kneel
knew|know
knitted|knit
knitting|knit
knobbed|knob
knobbing|knob
knotted|knot
knotting|knot
known|know
ko'd|ko
ko'ing|ko
ko's|ko
labelled|label
labelling|label
laden|lade
ladyfied|ladify
ladyfies|ladify
ladyfying|ladify
lagged|lag
lagging|lag
laid|lay
lain|lie
lallygagged|lallygag
lallygagging|lallygag
lammed|lam
lamming|lam
lapidified|lapidify
lapped|lap
lapping|lap
laurelled|laurel
laurelling|laurel
layed_for|lie_for
laying_for|lie_for
lays_for|lie_for
lay|lie
leant|lean
leapfrogged|leapfrog
leapfrogging|leapfrog
leapt|leap
learnt|learn
leaves_undone|leave_undone
leaving_undone|leave_undone
led|lead
left_undone|leave_undone
left|leave
lent|lend
letting|let
levelled|level
levelling|level
levied|levy
libelled|libel
libelling|libel
lignified|lignify
lipped|lip
lipping|lip
liquefied|liquify
liquefies|liquify
liquefy|liquify
liquified|liquify
lit|light
lobbed|lob
lobbied|lobby
lobbing|lob
logged|log
logging|log
looked_towards|look_towards
looking_towards|look_towards
looks_towards|look_towards
lopped|lop
lopping|lop
lost|lose
lotted|lot
lotting|lot
lugged|lug
lugging|lug
lullabied|lullaby
lying|lie
machine-gunned|machine-gun
machine-gunning|machine-gun
madded|mad
madding|mad
made|make
magnified|magnify
manned|man
manning|man
manumitted|manumit
manumitting|manumit
mapped|map
mapping|map
marcelled|marcel
marcelling|marcel
marred|mar
married|marry
marring|mar
marshalled|marshal
marshalling|marshal
marvelled|marvel
marvelling|marvel
matted|mat
matting|mat
meant|mean
medalled|medal
medalling|medal
metalled|metal
metalling|metal
metrified|metrify
met|meet
might|may
militated_against|militate_against
militates_against|militate_against
militating_against|militate_against
mimicked|mimic
mimicking|mimic
minified|minify
misapplied|misapply
misbecame|misbecome
miscarried|miscarry
misdealt|misdeal
misfitted|misfit
misfitting|misfit
misgave|misgive
misgiven|misgive
mishitting|mishit
mislaid|mislay
misled|mislead
mispled|misplead
misspelt|misspell
misspent|misspend
mistaken|mistake
mistook|mistake
misunderstood|misunderstand
mobbed|mob
mobbing|mob
modelled|model
modelling|model
modified|modify
mollified|mollify
molten|melt
mopped|mop
mopping|mop
mortified|mortify
mown|mow
mudded|mud
muddied|muddy
mudding|mud
mugged|mug
mugging|mug
multiplied|multiply
mummed|mum
mummified|mummify
mumming|mum
mutinied|mutiny
mystified|mystify
nabbed|nab
nabbing|nab
nagged|nag
nagging|nag
napped|nap
napping|nap
netted|net
netting|net
nibbed|nib
nibbing|nib
nickelled|nickel
nickelling|nickel
nid-nodded|nid-nod
nid-nodding|nid-nod
nidified|nidify
nigrified|nigrify
nipped|nip
nipping|nip
nitrified|nitrify
nodded|nod
nodding|nod
non-prossed|non-pros
non-prosses|non-pros
non-prossing|non-pros
nonplussed|nonplus
nonplusses|nonplus
nonplussing|nonplus
notified|notify
nullified|nullify
nutted|nut
nutting|nut
objectified|objectify
occupied|occupy
occurred|occur
occurring|occur
offsetting|offset
omitted|omit
omitting|omit
ossified|ossify
outbidden|outbid
outbidding|outbid
outbred|outbreed
outcried|outcry
outcropped|outcrop
outcropping|outcrop
outdid|outdo
outdone|outdo
outdrawn|outdraw
outdrew|outdraw
outfitted|outfit
outfitting|outfit
outfought|outfight
outgassed|outgas
outgasses|outgas
outgassing|outgas
outgeneralled|outgeneral
outgeneralling|outgeneral
outgone|outgo
outgrew|outgrow
outgrown|outgrow
outlaid|outlay
outmanned|outman
outmanning|outman
outputted|output
outputting|output
outran|outrun
outridden|outride
outrode|outride
outrunning|outrun
outshone|outshine
outshot|outshoot
outsold|outsell
outspanned|outspan
outspanning|outspan
outstood|outstand
outstripped|outstrip
outstripping|outstrip
outthought|outthink
outwent|outgo
outwitted|outwit
outwitting|outwit
outwore|outwear
outworn|outwear
overbidden|overbid
overbidding|overbid
overblew|overblow
overblown|overblow
overbore|overbear
overborne|overbear
overbuilt|overbuild
overcame|overcome
overcropped|overcrop
overcropping|overcrop
overdid|overdo
overdone|overdo
overdrawn|overdraw
overdrew|overdraw
overdriven|overdrive
overdrove|overdrive
overflew|overfly
overflown|overflow
overfly|overflow
overgrew|overgrow
overgrown|overgrow
overheard|overhear
overhung|overhang
overlaid|overlay
overlain|overlie
overlapped|overlap
overlapping|overlap
overlay|overlie
overlying|overlie
overmanned|overman
overmanning|overman
overpaid|overpay
overpast|overpass
overran|overrun
overridden|override
overrode|override
overrunning|overrun
oversaw|oversee
overseen|oversee
oversetting|overset
oversewn|oversew
overshot|overshoot
oversimplified|oversimplify
overslept|oversleep
oversold|oversell
overspent|overspend
overspilt|overspill
overstepped|overstep
overstepping|overstep
overtaken|overtake
overthrew|overthrow
overthrown|overthrow
overtook|overtake
overtopped|overtop
overtopping|overtop
overwound|overwind
overwritten|overwrite
overwrote|overwrite
pacified|pacify
padded|pad
padding|pad
paid|pay
palled|pal
palling|pal
palsied|palsy
pandied|pandy
panelled|panel
panelling|panel
panicked|panic
panicking|panic
panned|pan
panning|pan
parallelled|parallel
parallelling|parallel
parcelled|parcel
parcelling|parcel
parodied|parody
parried|parry
partaken|partake
partook|partake
pasquilled|pasquinade
pasquilling|pasquinade
pasquils|pasquinade
pasquil|pasquinade
patrolled|patrol
patrolling|patrol
patted|pat
patting|pat
pedalled|pedal
pedalling|pedal
pegged|peg
pegging|peg
pencilled|pencil
pencilling|pencil
penned|pen
penning|pen
pent|pen
pepped|pep
pepping|pep
permitted|permit
permitting|permit
personified|personify
petrified|petrify
petted|pet
pettifogged|pettifog
pettifogging|pettifog
petting|pet
phantasied|phantasy
photocopied|photocopy
photomapped|photomap
photomapping|photomap
photosetting|photoset
physicked|physic
physicking|physic
picnicked|picnic
picnicking|picnic
pigged|pig
pigging|pig
pilloried|pillory
pinch-hitting|pinch-hit
pinned|pin
pinning|pin
pipped|pip
pipping|pip
pistol-whipped|pistol-whip
pistol-whipping|pistol-whip
pistolled|pistol
pistolling|pistol
pitapatted|pitapat
pitapatting|pitapat
pitied|pity
pitted|pit
pitting|pit
planned|plan
planning|plan
platted|plat
platting|plat
played_a_part|play_a_part
playing_a_part|play_a_part
plays_a_part|play_a_part
pled|plead
plied|ply
plodded|plod
plodding|plod
plopped|plop
plopping|plop
plotted|plot
plotting|plot
plugged|plug
plugging|plug
podded|pod
podding|pod
pommelled|pommel
pommelling|pommel
popes|popes
popped|pop
popping|pop
potted|pot
potting|pot
preachified|preachify
precancelled|precancel
precancelling|precancel
preferred|prefer
preferring|prefer
preoccupied|preoccupy
prepaid|prepay
presignified|presignify
pretermitted|pretermit
pretermitting|pretermit
prettied|pretty
prettified|prettify
pried|pry
prigged|prig
prigging|prig
primmed|prim
primming|prim
prodded|prod
prodding|prod
programmed|program
programmes|program
programming|program
prologed|prologue
prologing|prologue
prologs|prologue
propelled|propel
propelling|propel
prophesied|prophesy
propped|prop
propping|prop
proven|prove
pubbed|pub
pubbing|pub
pugged|pug
pugging|pug
pummelled|pummel
pummelling|pummel
punned|pun
punning|pun
pupped|pup
pupping|pup
purified|purify
put-putted|put-put
put-putting|put-put
putrefied|putrefy
puttied|putty
putting|put
qualified|qualify
quantified|quantify
quarrelled|quarrel
quarrelling|quarrel
quarried|quarry
quartersawn|quartersaw
queried|query
quick-frozen|quick-freeze
quick-froze|quick-freeze
quickstepped|quickstep
quickstepping|quickstep
quipped|quip
quipping|quip
quitted|quit
quitting|quit
quizzed|quiz
quizzes|quiz
quizzing|quiz
ragged|rag
ragging|rag
rallied|rally
ramified|ramify
rammed|ram
ramming|ram
rang|ring
ran|run
rapped|rap
rappelled|rappel
rappelling|rappel
rapping|rap
rarefied|rarefy
ratified|ratify
ratted|rat
ratting|rat
ravelled|ravel
ravelling|ravel
razor-cutting|razor-cut
re-trodden|re-tread
re-trod|re-tread
rebelled|rebel
rebelling|rebel
rebuilt|rebuild
rebutted|rebut
rebutting|rebut
recapped|recap
recapping|recap
reclassified|reclassify
recommitted|recommit
recommitting|recommit
recopied|recopy
rectified|rectify
recurred|recur
recurring|recur
red-pencilled|red-pencil
red-pencilling|red-pencil
redded|red
redding|red
redd|red
redid|redo
redone|redo
red|red
referred|refer
referring|refer
refitted|refit
refitting|refit
reft|reave
refuelled|refuel
refuelling|refuel
regretted|regret
regretting|regret
reheard|rehear
reified|reify
relied|rely
remade|remake
remarried|remarry
remitted|remit
remitting|remit
rent|rend
repaid|repay
repelled|repel
repelling|repel
replevied|replevy
replied|reply
repotted|repot
repotting|repot
reran|rerun
rerunning|rerun
resat|resit
resetting|reset
resewn|resew
resitting|resit
retaken|retake
rethought|rethink
retold|retell
retook|retake
retransmitted|retransmit
retransmitting|retransmit
retried|retry
retrofitted|retrofit
retrofitting|retrofit
retted|ret
retting|ret
reunified|reunify
revelled|revel
revelling|revel
revetted|revet
revetting|revet
revivified|revivify
revved|rev
revving|rev
rewound|rewind
rewritten|rewrite
rewrote|rewrite
ribbed|rib
ribbing|rib
ricochetted|ricochet
ricochetting|ricochet
ridded|rid
ridden|ride
ridding|rid
rigged|rig
rigging|rig
rigidified|rigidify
rimmed|rim
rimming|rim
ripped|rip
ripping|rip
risen|rise
rivalled|rival
rivalling|rival
riven|rive
robbed|rob
robbing|rob
rode|ride
rose|rise
rotted|rot
rotting|rot
rough-dried|rough-dry
rough-hewn|rough-hew
rove|reeve
rowelled|rowel
rowelling|rowel
rubbed|rub
rubbing|rub
rung|ring
running|run
rutted|rut
rutting|rut
saccharified|saccharify
sagged|sag
sagging|sag
said|say
salaried|salary
salified|salify
sallied|sally
sanctified|sanctify
sandbagged|sandbag
sandbagging|sandbag
sang|sing
sank|sink
saponified|saponify
sapped|sap
sapping|sap
satisfied|satisfy
sat|sit
savvied|savvy
sawn|saw
saw|see
scagged|scag
scagging|scag
scanned|scan
scanning|scan
scarified|scarify
scarred|scar
scarring|scar
scatted|scat
scatting|scat
scorified|scorify
scragged|scrag
scragging|scrag
scrammed|scram
scramming|scram
scrapped|scrap
scrapping|scrap
scried|scry
scrubbed|scrub
scrubbing|scrub
scrummed|scrum
scrumming|scrum
scudded|scud
scudding|scud
scummed|scum
scumming|scum
scurried|scurry
seed|seed
seen|see
sent|send
setting|set
sewn|sew
shagged|shag
shagging|shag
shaken_hands|shake_hands
shaken|shake
shakes_hands|shake_hands
shaking_hands|shake_hands
shammed|sham
shamming|sham
sharecropped|sharecrop
sharecropping|sharecrop
shat|shit
shaven|shave
shedding|shed
shed|shed
shellacked|shellac
shellacking|shellac
shent|shend
shewn|shew
shied|shy
shikarred|shikar
shikarring|shikar
shillyshallied|shillyshally
shimmed|shim
shimmied|shimmy
shimming|shim
shinned|shin
shinning|shin
shipped|ship
shipping|ship
shitted|shit
shitting|shit
shod|shoe
shone|shine
shook_hands|shake_hands
shook|shake
shopped|shop
shopping|shop
shotgunned|shotgun
shotgunning|shotgun
shotted|shot
shotting|shot
shot|shoot
shovelled|shovel
shovelling|shovel
shown|show
shrank|shrink
shredded|shred
shredding|shred
shrink-wrapped|shrink-wrap
shrink-wrapping|shrink-wrap
shrivelled|shrivel
shrivelling|shrivel
shriven|shrive
shrove|shrive
shrugged|shrug
shrugging|shrug
shrunken|shrink
shrunk|shrink
shunned|shun
shunning|shun
shutting|shut
sicked|sic
sicking|sic
sideslipped|sideslip
sideslipping|sideslip
sidestepped|sidestep
sidestepping|sidestep
sightsaw|sightsee
sightseen|sightsee
signalled|signal
signalling|signal
signified|signify
silicified|silicify
simplified|simplify
singe|sing
singing|sing
single-stepped|single-step
single-stepping|single-step
sinned|sin
sinning|sin
sipped|sip
sipping|sip
sitting|sit
skellied|skelly
skenned|sken
skenning|sken
sketted|sket
sketting|sket
ski'd|ski
skidded|skid
skidding|skid
skimmed|skim
skimming|skim
skin-popped|skin-pop
skin-popping|skin-pop
skinned|skin
skinning|skin
skinny-dipped|skinny-dip
skinny-dipping|skinny-dip
skipped|skip
skipping|skip
skivvied|skivvy
skydove|skydive
slabbed|slab
slabbing|slab
slagged|slag
slagging|slag
slain|slay
slammed|slam
slamming|slam
slapped|slap
slapping|slap
slatted|slat
slatting|slat
sledding|sled
slept|sleep
slew|slay
slidden|slide
slid|slide
slimming|slim
slipped|slip
slipping|slip
slitting|slit
slogged|slog
slogging|slog
slopped|slop
slopping|slop
slotted|slot
slotting|slot
slugged|slug
slugging|slug
slummed|slum
slumming|slum
slung|sling
slunk|slink
slurred|slur
slurring|slur
smelt|smell
smitten|smite
smit|smite
smote|smite
smutted|smut
smutting|smut
snagged|snag
snagging|snag
snapped|snap
snapping|snap
snedded|sned
snedding|sned
snipped|snip
snipping|snip
snivelled|snivel
snivelling|snivel
snogged|snog
snogging|snog
snubbed|snub
snubbing|snub
snuck|sneak
snugged|snug
snugging|snug
sobbed|sob
sobbing|sob
sodded|sod
sodding|sod
soft-pedalled|soft-pedal
soft-pedalling|soft-pedal
sold|sell
solemnified|solemnify
solidified|solidify
soothsaid|soothsay
sopped|sop
sopping|sop
sought|seek
sown|sow
spagged|spag
spagging|spag
spancelled|spancel
spancelling|spancel
spanned|span
spanning|span
sparred|spar
sparring|spar
spatted|spat
spatting|spat
spat|spit
specified|specify
sped|speed
speechified|speechify
spellbound|spellbind
spelt|spell
spent|spend
spied|spy
spilt|spill
spin-dried|spin-dry
spinning|spin
spiralled|spiral
spiralling|spiral
spitted|spit
spitting|spit
splitting|split
spoilt|spoil
spoken|speak
spoke|speak
spoon-fed|spoon-feed
spotlit|spotlight
spotted|spot
spotting|spot
sprang|spring
sprigged|sprig
sprigging|sprig
sprung|spring
spudded|spud
spudding|spud
spun|spin
spurred|spur
spurring|spur
squatted|squat
squatting|squat
squibbed|squib
squibbing|squib
squidded|squid
squidding|squid
squilgee|squeegee
stabbed|stab
stabbing|stab
stall-fed|stall-feed
stank|stink
starred|star
starring|star
steadied|steady
stellified|stellify
stemmed|stem
stemming|stem
stems_from|stem_from
stencilled|stencil
stencilling|stencil
stepped|step
stepping|step
stetted|stet
stetting|stet
stied|sty
stilettoeing|stiletto
stirred|stir
stirring|stir
stolen|steal
stole|steal
stood|stand
stopped|stop
stopping|stop
storied|story
stotted|stot
stotting|stot
stove|stave
strapped|strap
strapping|strap
stratified|stratify
strewn|strew
stricken|strike
stridden|stride
stripped|strip
stripping|strip
striven|strive
strode|stride
stropped|strop
stropping|strop
strove|strive
strown|strow
struck|strike
strummed|strum
strumming|strum
strung|string
strutted|strut
strutting|strut
stubbed|stub
stubbing|stub
stuck|stick
studded|stud
studding|stud
studied|study
stultified|stultify
stummed|stum
stumming|stum
stung|sting
stunk|stink
stunned|stun
stunning|stun
stupefied|stupefy
stymying|stymie
subbed|sub
subbing|sub
subjectified|subjectify
subletting|sublet
submitted|submit
submitting|submit
subtotalled|subtotal
subtotalling|subtotal
sullied|sully
sulphuretted|sulphuret
sulphuretting|sulphuret
summed|sum
summing|sum
sung|sing
sunken|sink
sunk|sink
sunned|sun
sunning|sun
supped|sup
supping|sup
supplied|supply
swabbed|swab
swabbing|swab
swagged|swag
swagging|swag
swam|swim
swapped|swap
swapping|swap
swatted|swat
swatting|swat
swept|sweep
swigged|swig
swigging|swig
swimming|swim
swivelled|swivel
swivelling|swivel
swollen|swell
swopped|swap
swopping|swap
swops|swap
swore|swear
sworn|swear
swotted|swot
swotting|swot
swum|swim
swung|swing
syllabified|syllabify
symbolled|symbol
symbolling|symbol
tabbed|tab
tabbing|tab
tagged|tag
tagging|tag
taken_a_side|take_a_side
taken_pains|take_pains
taken_steps|take_steps
taken|take
takes_a_side|take_a_side
takes_pains|take_pains
takes_steps|take_steps
taking_a_side|take_a_side
taking_pains|take_pains
taking_steps|take_steps
talcked|talc
talcking|talc
tallied|tally
tally-ho'd|tally-ho
tammied|tammy
tanned|tan
tanning|tan
tapped|tap
tapping|tap
tarred|tar
tarried|tarry
tarring|tar
tasselled|tassel
tasselling|tassel
tatted|tat
tatting|tat
taught|teach
taxis|taxis
taxying|taxi
teaselled|teasel
teaselling|teasel
tedded|ted
tedding|ted
tepefied|tepefy
terrified|terrify
testes|testes
testified|testify
thinking_the_world_of|think_the_world_of
thinks_the_world_of|think_the_world_of
thinned|thin
thinning|thin
thought_the_world_of|think_the_world_of
thought|think
threw_out|throw_out
threw|throw
thriven|thrive
throbbed|throb
throbbing|throb
throve|thrive
throwing_out|throw_out
thrown_out|throw_out
thrown|throw
throws_out|throw_out
thrummed|thrum
thrumming|thrum
thudded|thud
thudding|thud
thwapping|thwap
tidied|tidy
tinned|tin
tinning|tin
tinselled|tinsel
tinselling|tinsel
tipped|tip
tipping|tip
tittupped|tittup
tittupping|tittup
toadied|toady
togged|tog
togging|tog
told|tell
took_a_side|take_a_side
took_pains|take_pains
took_steps|take_steps
took|take
topped|top
topping|top
tore|tear
torn|tear
torrefied|torrefy
torrify|torrefy
totalled|total
totalling|total
totted|tot
totting|tot
towelled|towel
towelling|towel
trafficked|traffic
trafficking|traffic
trameled|trammel
trameling|trammel
tramelled|trammel
tramelling|trammel
tramels|trammel
trammed|tram
tramming|tram
transferred|transfer
transferring|transfer
transfixt|transfix
transhipped|tranship
transhipping|tranship
tranship|transship
transmitted|transmit
transmitting|transmit
transmogrified|transmogrify
transshipped|transship
transshipping|transship
trapanned|trapan
trapanning|trapan
trapped|trap
trapping|trap
travelled|travel
travelling|travel
travestied|travesty
trekked|trek
trekking|trek
trepanned|trepan
trepanning|trepan
tried|try
trigged|trig
trigging|trig
trimmed|trim
trimming|trim
tripped|trip
tripping|trip
trodden|tread
trod|tread
trogged|trog
trogging|trog
trotted|trot
trotting|trot
trowelled|trowel
trowelling|trowel
tugged|tug
tugging|tug
tumefied|tumefy
tunned|tun
tunnelled|tunnel
tunnelling|tunnel
tunning|tun
tupped|tup
tupping|tup
tut-tutted|tut-tut
tut-tutting|tut-tut
twigged|twig
twigging|twig
twinned|twin
twinning|twin
twitted|twit
twitting|twit
tying|tie
typesetting|typeset
typewritten|typewrite
typewrote|typewrite
typified|typify
uglified|uglify
unbarred|unbar
unbarring|unbar
unbent|unbend
unbound|unbind
uncapped|uncap
uncapping|uncap
unclad|unclothe
unclogged|unclog
unclogging|unclog
underbidding|underbid
underbought|underbuy
undercutting|undercut
underfed|underfeed
undergirt|undergird
undergone|undergo
underlaid|underlay
underlain|underlie
underlay|underlie
underletting|underlet
underlying|underlie
underpaid|underpay
underpinned|underpin
underpinning|underpin
underpropped|underprop
underpropping|underprop
undersetting|underset
undershot|undershoot
undersold|undersell
understood|understand
understudied|understudy
undertaken|undertake
undertook|undertake
underwent|undergo
underwritten|underwrite
underwrote|underwrite
undid|undo
undone|undo
unfitted|unfit
unfitting|unfit
unfrozen|unfreeze
unfroze|unfreeze
unified|unify
unkennelled|unkennel
unkennelling|unkennel
unknitted|unknit
unknitting|unknit
unlaid|unlay
unlearnt|unlearn
unmade|unmake
unmanned|unman
unmanning|unman
unpegged|unpeg
unpegging|unpeg
unpinned|unpin
unpinning|unpin
unplugged|unplug
unplugging|unplug
unravelled|unravel
unravelling|unravel
unrigged|unrig
unrigging|unrig
unripped|unrip
unripping|unrip
unrove|unreeve
unsaid|unsay
unshipped|unship
unshipping|unship
unslung|unsling
unsnapped|unsnap
unsnapping|unsnap
unspoken|unspeak
unspoke|unspeak
unsteadied|unsteady
unstepped|unstep
unstepping|unstep
unstopped|unstop
unstopping|unstop
unstrung|unstring
unstuck|unstick
unswore|unswear
unsworn|unswear
untaught|unteach
unthought|unthink
untidied|untidy
untrodden|untread
untrod|untread
untying|untie
unwound|unwind
unwrapped|unwrap
unwrapping|unwrap
unzipped|unzip
unzipping|unzip
upbuilt|upbuild
upheld|uphold
uphove|upheave
upped|up
uppercutting|uppercut
upping|up
uprisen|uprise
uprose|uprise
upsetting|upset
upsprang|upspring
upsprung|upspring
upswept|upsweep
upswollen|upswell
upswung|upswing
vagged|vag
vagging|vag
varied|vary
vatted|vat
vatting|vat
verbified|verbify
verified|verify
versified|versify
vetted|vet
vetting|vet
victualled|victual
victualling|victual
vilified|vilify
vitrified|vitrify
vitriolled|vitriol
vitriolling|vitriol
vivified|vivify
vying|vie
wadded|wad
waddied|waddy
wadding|wad
wadsetted|wadset
wadsetting|wadset
wagged|wag
wagging|wag
wanned|wan
wanning|wan
warred|war
warring|war
was|be
water-ski'd|water-ski
waylaid|waylay
wearied|weary
weatherstripped|weatherstrip
weatherstripping|weatherstrip
webbed|web
webbing|web
wedded|wed
wedding|wed
weed|weed
went_deep|go_deep
went|go
wept|weep
were|be
wetted|wet
wetting|wet
whammed|wham
whamming|wham
whapped|whap
whapping|whap
whetted|whet
whetting|whet
whinnied|whinny
whipped|whip
whipping|whip
whipsawn|whipsaw
whirred|whir
whirring|whir
whistle-stopped|whistle-stop
whistle-stopping|whistle-stop
whizzed|whiz
whizzes|whiz
whizzing|whiz
whopped|whop
whopping|whop
wigged|wig
wigging|wig
wigwagged|wigwag
wigwagging|wigwag
wildcatted|wildcat
wildcatting|wildcat
window-shopped|window-shop
window-shopping|window-shop
winning|win
winterfed|winterfeed
wiredrawn|wiredraw
wiredrew|wiredraw
withdrawn|withdraw
withdrew|withdraw
withheld|withhold
withstood|withstand
woken|wake
woke|wake
wonned|won
wonning|won
won|win
wore|wear
worn|wear
worried|worry
worshipped|worship
worshipping|worship
wound|wind
woven|weave
wove|weave
wrapped|wrap
wrapping|wrap
wried|wry
written|write
wrote|write
wrought|work
wrung|wring
yakked|yak
yakking|yak
yapped|yap
yapping|yap
ycleped|clepe
yclept|clepe
yenned|yen
yenning|yen
yodelled|yodel
yodelling|yodel
zapped|zap
zapping|zap
zigzagged|zigzag
zigzagging|zigzag
zipped|zip
zipping|zip